//
// PCILeech FPGA.
//
// PCIe BAR PIO controller.
//
// The PCILeech BAR PIO controller allows for easy user-implementation on top
// of the PCILeech AXIS128 PCIe TLP streaming interface.
// The controller consists of a read engine and a write engine and pluggable
// user-implemented PCIe BAR implementations (found at bottom of the file).
//
// Considerations:
// - The core handles 1 DWORD read + 1 DWORD write per CLK max. If a lot of
//   data is written / read from the TLP streaming interface the core may
//   drop packet silently.
// - The core reads 1 DWORD of data (without byte enable) per CLK.
// - The core writes 1 DWORD of data (with byte enable) per CLK.
// - All user-implemented cores must have the same latency in CLKs for the
//   returned read data or else undefined behavior will take place.
// - 32-bit addresses are passed for read/writes. Larger BARs than 4GB are
//   not supported due to addressing constraints. Lower bits (LSBs) are the
//   BAR offset, Higher bits (MSBs) are the 32-bit base address of the BAR.
// - DO NOT edit read/write engines.
// - DO edit pcileech_tlps128_bar_controller (to swap bar implementations).
// - DO edit the bar implementations (at bottom of the file, if neccessary).
//
// Example implementations exists below, swap out any of the example cores
// against a core of your use case, or modify existing cores.
// Following test cores exist (see below in this file):
// - pcileech_bar_impl_zerowrite4k = zero-initialized read/write BAR.
//     It's possible to modify contents by use of .coe file.
// - pcileech_bar_impl_loopaddr = test core that loops back the 32-bit
//     address of the current read. Does not support writes.
// - pcileech_bar_impl_none = core without any reply.
// 
// (c) Ulf Frisk, 2024
// Author: Ulf Frisk, pcileech@frizk.net
//

`timescale 1ns / 1ps
`include "pcileech_header.svh"

module pcileech_tlps128_bar_controller(
    input                   rst,
    input                   clk,
    input                   bar_en,
    input [15:0]            pcie_id,
    IfAXIS128.sink_lite     tlps_in,
    IfAXIS128.source        tlps_out,
    output                  int_enable,
    input                   msix_vaild,
    output                  msix_send_done,
    output [31:0]           msix_address,
    output [31:0]           msix_vector,
    input [31:0]            base_address_register,
    input [31:0]            base_address_register_1,
    input [31:0]            base_address_register_2,
    input [31:0]            base_address_register_3,
    input [31:0]            base_address_register_4,
    input [31:0]            base_address_register_5
);
    
    // ------------------------------------------------------------------------
    // 1: TLP RECEIVE:
    // Receive incoming BAR requests from the TLP stream:
    // send them onwards to read and write FIFOs
    // ------------------------------------------------------------------------
    wire in_is_wr_ready;
    bit  in_is_wr_last;
    wire in_is_first    = tlps_in.tuser[0];
    wire in_is_bar      = bar_en && (tlps_in.tuser[8:2] != 0);
    wire in_is_rd       = (in_is_first && tlps_in.tlast && ((tlps_in.tdata[31:25] == 7'b0000000) || (tlps_in.tdata[31:25] == 7'b0010000) || (tlps_in.tdata[31:24] == 8'b00000010)));
    wire in_is_wr       = in_is_wr_last || (in_is_first && in_is_wr_ready && ((tlps_in.tdata[31:25] == 7'b0100000) || (tlps_in.tdata[31:25] == 7'b0110000) || (tlps_in.tdata[31:24] == 8'b01000010)));
    
    always @ ( posedge clk )
        if ( rst ) begin
            in_is_wr_last <= 0;
        end
        else if ( tlps_in.tvalid ) begin
            in_is_wr_last <= !tlps_in.tlast && in_is_wr;
        end
    
    wire [6:0]  wr_bar;
    wire [31:0] wr_addr;
    wire [3:0]  wr_be;
    wire [31:0] wr_data;
    wire        wr_valid;
    wire [87:0] rd_req_ctx;
    wire [6:0]  rd_req_bar;
    wire [31:0] rd_req_addr;
    wire [3:0]  rd_req_be;
    wire        rd_req_valid;
    wire [87:0] rd_rsp_ctx;
    wire [31:0] rd_rsp_data;
    wire        rd_rsp_valid;
        
    pcileech_tlps128_bar_rdengine i_pcileech_tlps128_bar_rdengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .pcie_id        ( pcie_id                       ),
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_rd ),
        .tlps_out       ( tlps_out                      ),
        // BAR reads:
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_bar     ( rd_req_bar                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_be      ( rd_req_be                     ),
        .rd_req_valid   ( rd_req_valid                  ),
        .rd_rsp_ctx     ( rd_rsp_ctx                    ),
        .rd_rsp_data    ( rd_rsp_data                   ),
        .rd_rsp_valid   ( rd_rsp_valid                  )
    );

    pcileech_tlps128_bar_wrengine i_pcileech_tlps128_bar_wrengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_wr ),
        .tlps_in_ready  ( in_is_wr_ready                ),
        // outgoing BAR writes:
        .wr_bar         ( wr_bar                        ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid                      )
    );
    
    wire [87:0] bar_rsp_ctx[7];
    wire [31:0] bar_rsp_data[7];
    wire        bar_rsp_valid[7];
    
    assign rd_rsp_ctx = bar_rsp_valid[0] ? bar_rsp_ctx[0] :
                        bar_rsp_valid[1] ? bar_rsp_ctx[1] :
                        bar_rsp_valid[2] ? bar_rsp_ctx[2] :
                        bar_rsp_valid[3] ? bar_rsp_ctx[3] :
                        bar_rsp_valid[4] ? bar_rsp_ctx[4] :
                        bar_rsp_valid[5] ? bar_rsp_ctx[5] :
                        bar_rsp_valid[6] ? bar_rsp_ctx[6] : 0;
    assign rd_rsp_data = bar_rsp_valid[0] ? bar_rsp_data[0] :
                        bar_rsp_valid[1] ? bar_rsp_data[1] :
                        bar_rsp_valid[2] ? bar_rsp_data[2] :
                        bar_rsp_valid[3] ? bar_rsp_data[3] :
                        bar_rsp_valid[4] ? bar_rsp_data[4] :
                        bar_rsp_valid[5] ? bar_rsp_data[5] :
                        bar_rsp_valid[6] ? bar_rsp_data[6] : 0;
    assign rd_rsp_valid = bar_rsp_valid[0] || bar_rsp_valid[1] || bar_rsp_valid[2] || bar_rsp_valid[3] || bar_rsp_valid[4] || bar_rsp_valid[5] || bar_rsp_valid[6];
    
    
    
    // 这是一个模拟
    assign int_enable = 1;
    
    pcileech_bar_impl_none i_bar0(
        .rst                   ( rst                           ),
        .clk                   ( clk                           ),
        .wr_addr               ( wr_addr                       ),
        .wr_be                 ( wr_be                         ),
        .wr_data               ( wr_data                       ),
        .wr_valid              ( wr_valid && wr_bar[0]         ),
        .rd_req_ctx            ( rd_req_ctx                    ),
        .rd_req_addr           ( rd_req_addr                   ),
        .rd_req_valid          ( rd_req_valid && rd_req_bar[0] ),
        .rd_rsp_ctx            ( bar_rsp_ctx[0]                ),
        .rd_rsp_data           ( bar_rsp_data[0]               ),
        .rd_rsp_valid          ( bar_rsp_valid[0]              )
    );
    
    pcileech_bar_impl_none i_bar1(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[1]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[1] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[1]                ),
        .rd_rsp_data    ( bar_rsp_data[1]               ),
        .rd_rsp_valid   ( bar_rsp_valid[1]              )
    );
    
    pcileech_bar_impl_bar2 i_bar2(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[2]         ),
        .base_address_register (base_address_register_2 ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[2] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[2]                ),
        .rd_rsp_data    ( bar_rsp_data[2]               ),
        .rd_rsp_valid   ( bar_rsp_valid[2]              )
    );
    
    pcileech_bar_impl_none i_bar3(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[3]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[3] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[3]                ),
        .rd_rsp_data    ( bar_rsp_data[3]               ),
        .rd_rsp_valid   ( bar_rsp_valid[3]              )
    );
    
    pcileech_bar_impl_bar4 i_bar4(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[4]         ),
        .base_address_register (base_address_register_4 ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[4] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[4]                ),
        .rd_rsp_data    ( bar_rsp_data[4]               ),
        .rd_rsp_valid   ( bar_rsp_valid[4]              )
    );
    
    pcileech_bar_impl_none i_bar5(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[5]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[5] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[5]                ),
        .rd_rsp_data    ( bar_rsp_data[5]               ),
        .rd_rsp_valid   ( bar_rsp_valid[5]              )
    );
    
    pcileech_bar_impl_none i_bar6_optrom(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[6]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[6] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[6]                ),
        .rd_rsp_data    ( bar_rsp_data[6]               ),
        .rd_rsp_valid   ( bar_rsp_valid[6]              )
    );


endmodule



// ------------------------------------------------------------------------
// BAR WRITE ENGINE:
// Receives BAR WRITE TLPs and output BAR WRITE requests.
// Holds a 2048-byte buffer.
// Input flow rate is 16bytes/CLK (max).
// Output flow rate is 4bytes/CLK.
// If write engine overflows incoming TLP is completely discarded silently.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_wrengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    output                  tlps_in_ready,
    // outgoing BAR writes:
    output bit [6:0]        wr_bar,
    output bit [31:0]       wr_addr,
    output bit [3:0]        wr_be,
    output bit [31:0]       wr_data,
    output bit              wr_valid
);

    wire            f_rd_en;
    wire [127:0]    f_tdata;
    wire [3:0]      f_tkeepdw;
    wire [8:0]      f_tuser;
    wire            f_tvalid;
    
    bit [127:0]     tdata;
    bit [3:0]       tkeepdw;
    bit             tlast;
    
    bit [3:0]       be_first;
    bit [3:0]       be_last;
    bit             first_dw;
    bit [31:0]      addr;

    fifo_141_141_clk1_bar_wr i_fifo_141_141_clk1_bar_wr(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( {tlps_in.tuser[8:0], tlps_in.tkeepdw, tlps_in.tdata} ),
        .full           (                               ),
        .prog_empty     ( tlps_in_ready                 ),
        .rd_en          ( f_rd_en                       ),
        .dout           ( {f_tuser, f_tkeepdw, f_tdata} ),    
        .empty          (                               ),
        .valid          ( f_tvalid                      )
    );
    
    // STATE MACHINE:
    `define S_ENGINE_IDLE        3'h0
    `define S_ENGINE_FIRST       3'h1
    `define S_ENGINE_4DW_REQDATA 3'h2
    `define S_ENGINE_TX0         3'h4
    `define S_ENGINE_TX1         3'h5
    `define S_ENGINE_TX2         3'h6
    `define S_ENGINE_TX3         3'h7
    (* KEEP = "TRUE" *) bit [3:0] state = `S_ENGINE_IDLE;
    
    assign f_rd_en = (state == `S_ENGINE_IDLE) ||
                     (state == `S_ENGINE_4DW_REQDATA) ||
                     (state == `S_ENGINE_TX3) ||
                     ((state == `S_ENGINE_TX2 && !tkeepdw[3])) ||
                     ((state == `S_ENGINE_TX1 && !tkeepdw[2])) ||
                     ((state == `S_ENGINE_TX0 && !f_tkeepdw[1]));

    always @ ( posedge clk ) begin
        wr_addr     <= addr;
        wr_valid    <= ((state == `S_ENGINE_TX0) && f_tvalid) || (state == `S_ENGINE_TX1) || (state == `S_ENGINE_TX2) || (state == `S_ENGINE_TX3);
        
    end

    always @ ( posedge clk )
        if ( rst ) begin
            state <= `S_ENGINE_IDLE;
        end
        else case ( state )
            `S_ENGINE_IDLE: begin
                state   <= `S_ENGINE_FIRST;
            end
            `S_ENGINE_FIRST: begin
                if ( f_tvalid && f_tuser[0] ) begin
                    wr_bar      <= f_tuser[8:2];
                    tdata       <= f_tdata;
                    tkeepdw     <= f_tkeepdw;
                    tlast       <= f_tuser[1];
                    first_dw    <= 1;
                    be_first    <= f_tdata[35:32];
                    be_last     <= f_tdata[39:36];
                    if ( f_tdata[31:29] == 8'b010 ) begin       // 3 DW header, with data
                        addr    <= { f_tdata[95:66], 2'b00 };
                        state   <= `S_ENGINE_TX3;
                    end
                    else if ( f_tdata[31:29] == 8'b011 ) begin  // 4 DW header, with data
                        addr    <= { f_tdata[127:98], 2'b00 };
                        state   <= `S_ENGINE_4DW_REQDATA;
                    end 
                end
                else begin
                    state   <= `S_ENGINE_IDLE;
                end
            end 
            `S_ENGINE_4DW_REQDATA: begin
                state   <= `S_ENGINE_TX0;
            end
            `S_ENGINE_TX0: begin
                tdata       <= f_tdata;
                tkeepdw     <= f_tkeepdw;
                tlast       <= f_tuser[1];
                addr        <= addr + 4;
                wr_data     <= { f_tdata[0+00+:8], f_tdata[0+08+:8], f_tdata[0+16+:8], f_tdata[0+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (f_tkeepdw[1] ? 4'hf : be_last);
                state       <= f_tvalid ? (f_tkeepdw[1] ? `S_ENGINE_TX1 : `S_ENGINE_FIRST) : `S_ENGINE_IDLE;
            end
            `S_ENGINE_TX1: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[32+00+:8], tdata[32+08+:8], tdata[32+16+:8], tdata[32+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[2] ? 4'hf : be_last);
                state       <= tkeepdw[2] ? `S_ENGINE_TX2 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX2: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[64+00+:8], tdata[64+08+:8], tdata[64+16+:8], tdata[64+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[3] ? 4'hf : be_last);
                state       <= tkeepdw[3] ? `S_ENGINE_TX3 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX3: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[96+00+:8], tdata[96+08+:8], tdata[96+16+:8], tdata[96+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (!tlast ? 4'hf : be_last);
                state       <= !tlast ? `S_ENGINE_TX0 : `S_ENGINE_FIRST;
            end
        endcase

endmodule




// ------------------------------------------------------------------------
// BAR READ ENGINE:
// Receives BAR READ TLPs and output BAR READ requests.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_rdengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    input [15:0]            pcie_id,
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    IfAXIS128.source        tlps_out,
    // BAR reads:
    output [87:0]           rd_req_ctx,
    output [6:0]            rd_req_bar,
    output [31:0]           rd_req_addr,
    output                  rd_req_valid,
    output [3:0]            rd_req_be,        
    input  [87:0]           rd_rsp_ctx,
    input  [31:0]           rd_rsp_data,
    input                   rd_rsp_valid
);
    // ------------------------------------------------------------------------
    // 1: PROCESS AND QUEUE INCOMING READ TLPs:
    // ------------------------------------------------------------------------
    wire [10:0] rd1_in_dwlen    = (tlps_in.tdata[9:0] == 0) ? 11'd1024 : {1'b0, tlps_in.tdata[9:0]};
    wire [6:0]  rd1_in_bar      = tlps_in.tuser[8:2];
    wire [15:0] rd1_in_reqid    = tlps_in.tdata[63:48];
    wire [7:0]  rd1_in_tag      = tlps_in.tdata[47:40];
    wire [31:0] rd1_in_addr     = { ((tlps_in.tdata[31:29] == 3'b000) ? tlps_in.tdata[95:66] : tlps_in.tdata[127:98]), 2'b00 };
    wire [3:0]  rd1_in_be       = tlps_in.tdata[35:32];
    wire [73:0] rd1_in_data;
    assign rd1_in_data[73:63]   = rd1_in_dwlen;
    assign rd1_in_data[62:56]   = rd1_in_bar;   
    assign rd1_in_data[55:48]   = rd1_in_tag;
    assign rd1_in_data[47:32]   = rd1_in_reqid;
    assign rd1_in_data[31:0]    = rd1_in_addr;

    
    wire [3:0]  rd1_out_be;
    wire        rd1_out_be_valid;
    wire        rd1_out_rden;
    wire [73:0] rd1_out_data;
    wire        rd1_out_valid;
    
    fifo_74_74_clk1_bar_rd1 i_fifo_74_74_clk1_bar_rd1(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( rd1_in_data                   ),
        .full           (                               ),
        .rd_en          ( rd1_out_rden                  ),
        .dout           ( rd1_out_data                  ),    
        .empty          (                               ),
        .valid          ( rd1_out_valid                 )
    );
    fifo_4_4_clk1_bar_rd1 i_fifo_4_4_clk1_bar_rd1 (
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( rd1_in_be                     ),
        .full           (                               ),
        .rd_en          ( rd1_out_rden                  ),
        .dout           ( rd1_out_be                    ),
        .empty          (                               ),
        .valid          ( rd1_out_be_valid              )

    );
    
    // ------------------------------------------------------------------------
    // 2: PROCESS AND SPLIT READ TLPs INTO RESPONSE TLP READ REQUESTS AND QUEUE:
    //    (READ REQUESTS LARGER THAN 128-BYTES WILL BE SPLIT INTO MULTIPLE).
    // ------------------------------------------------------------------------
    
    wire [10:0] rd1_out_dwlen       = rd1_out_data[73:63];
    wire [4:0]  rd1_out_dwlen5      = rd1_out_data[67:63];
    wire [4:0]  rd1_out_addr5       = rd1_out_data[6:2];
    
    // 1st "instant" packet:
    wire [4:0]  rd2_pkt1_dwlen_pre  = ((rd1_out_addr5 + rd1_out_dwlen5 > 6'h20) || ((rd1_out_addr5 != 0) && (rd1_out_dwlen5 == 0))) ? (6'h20 - rd1_out_addr5) : rd1_out_dwlen5;
    wire [5:0]  rd2_pkt1_dwlen      = (rd2_pkt1_dwlen_pre == 0) ? 6'h20 : rd2_pkt1_dwlen_pre;
    wire [10:0] rd2_pkt1_dwlen_next = rd1_out_dwlen - rd2_pkt1_dwlen;
    wire        rd2_pkt1_large      = (rd1_out_dwlen > 32) || (rd1_out_dwlen != rd2_pkt1_dwlen);
    wire        rd2_pkt1_tiny       = (rd1_out_dwlen == 1);
    wire [11:0] rd2_pkt1_bc         = rd1_out_dwlen << 2;
    wire [85:0] rd2_pkt1;
    assign      rd2_pkt1[85:74]     = rd2_pkt1_bc;
    assign      rd2_pkt1[73:63]     = rd2_pkt1_dwlen;
    assign      rd2_pkt1[62:0]      = rd1_out_data[62:0];
    
    // Nth packet (if split should take place):
    bit  [10:0] rd2_total_dwlen;
    wire [10:0] rd2_total_dwlen_next = rd2_total_dwlen - 11'h20;
    
    bit  [85:0] rd2_pkt2;
    wire [10:0] rd2_pkt2_dwlen = rd2_pkt2[73:63];
    wire        rd2_pkt2_large = (rd2_total_dwlen > 11'h20);
    
    wire        rd2_out_rden;
    
    // STATE MACHINE:
    `define S2_ENGINE_REQDATA     1'h0
    `define S2_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state2 = `S2_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            state2 <= `S2_ENGINE_REQDATA;
        end
        else case ( state2 )
            `S2_ENGINE_REQDATA: begin
                if ( rd1_out_valid && rd2_pkt1_large ) begin
                    rd2_total_dwlen <= rd2_pkt1_dwlen_next;                             // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_pkt1_dwlen_next << 2;                        // byte-count
                    rd2_pkt2[73:63] <= (rd2_pkt1_dwlen_next > 11'h20) ? 11'h20 : rd2_pkt1_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd1_out_data[62:12];                             // various data
                    rd2_pkt2[11:0]  <= rd1_out_data[11:0] + (rd2_pkt1_dwlen << 2);      // base address (within 4k page)
                    state2 <= `S2_ENGINE_PROCESSING;
                end
            end
            `S2_ENGINE_PROCESSING: begin
                if ( rd2_out_rden ) begin
                    rd2_total_dwlen <= rd2_total_dwlen_next;                                // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_total_dwlen_next << 2;                           // byte-count
                    rd2_pkt2[73:63] <= (rd2_total_dwlen_next > 11'h20) ? 11'h20 : rd2_total_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd2_pkt2[62:12];                                     // various data
                    rd2_pkt2[11:0]  <= rd2_pkt2[11:0] + (rd2_pkt2_dwlen << 2);              // base address (within 4k page)
                    if ( !rd2_pkt2_large ) begin
                        state2 <= `S2_ENGINE_REQDATA;
                    end
                end
            end
        endcase
    
    assign rd1_out_rden = rd2_out_rden && (((state2 == `S2_ENGINE_REQDATA) && (!rd1_out_valid || rd2_pkt1_tiny)) || ((state2 == `S2_ENGINE_PROCESSING) && !rd2_pkt2_large));

    wire [85:0] rd2_in_data  = (state2 == `S2_ENGINE_REQDATA) ? rd2_pkt1 : rd2_pkt2;
    wire        rd2_in_valid = rd1_out_valid || ((state2 == `S2_ENGINE_PROCESSING) && rd2_out_rden);
    wire [3:0]  rd2_in_be       = rd1_out_be;
    wire        rd2_in_be_valid = rd1_out_valid;

    bit  [85:0] rd2_out_data;
    bit         rd2_out_valid;
    bit  [3:0]  rd2_out_be;
    bit         rd2_out_be_valid;
    always @ ( posedge clk ) begin
        rd2_out_data    <= rd2_in_valid ? rd2_in_data : rd2_out_data;
        rd2_out_valid   <= rd2_in_valid && !rst;
        rd2_out_be       <= rd2_in_be_valid ? rd2_in_be : rd2_out_data;
        rd2_out_be_valid <= rd2_in_be_valid && !rst;  
    end

    // ------------------------------------------------------------------------
    // 3: PROCESS EACH READ REQUEST PACKAGE PER INDIVIDUAL 32-bit READ DWORDS:
    // ------------------------------------------------------------------------

    wire [4:0]  rd2_out_dwlen   = rd2_out_data[67:63];
    wire        rd2_out_last    = (rd2_out_dwlen == 1);
    wire [9:0]  rd2_out_dwaddr  = rd2_out_data[11:2];
    
    wire        rd3_enable;
    
    bit [3:0]   rd3_process_be;
    bit         rd3_process_valid;
    bit         rd3_process_first;
    bit         rd3_process_last;
    bit [4:0]   rd3_process_dwlen;
    bit [9:0]   rd3_process_dwaddr;
    bit [85:0]  rd3_process_data;
    wire        rd3_process_next_last = (rd3_process_dwlen == 2);
    wire        rd3_process_nextnext_last = (rd3_process_dwlen <= 3);
    assign rd_req_be    = rd3_process_be;
    assign rd_req_ctx   = { rd3_process_first, rd3_process_last, rd3_process_data };
    assign rd_req_bar   = rd3_process_data[62:56];
    assign rd_req_addr  = { rd3_process_data[31:12], rd3_process_dwaddr, 2'b00 };
    assign rd_req_valid = rd3_process_valid;
    
    // STATE MACHINE:
    `define S3_ENGINE_REQDATA     1'h0
    `define S3_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state3 = `S3_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            rd3_process_valid   <= 1'b0;
            state3              <= `S3_ENGINE_REQDATA;
        end
        else case ( state3 )
            `S3_ENGINE_REQDATA: begin
                if ( rd2_out_valid ) begin
                    rd3_process_valid       <= 1'b1;
                    rd3_process_first       <= 1'b1;                    // FIRST
                    rd3_process_last        <= rd2_out_last;            // LAST (low 5 bits of dwlen == 1, [max pktlen = 0x20))
                    rd3_process_dwlen       <= rd2_out_dwlen;           // PKT LENGTH IN DW
                    rd3_process_dwaddr      <= rd2_out_dwaddr;          // DWADDR OF THIS DWORD
                    rd3_process_data[85:0]  <= rd2_out_data[85:0];      // FORWARD / SAVE DATA
                    if ( rd2_out_be_valid ) begin
                        rd3_process_be <= rd2_out_be;
                    end else begin
                        rd3_process_be <= 4'hf;
                    end
                    if ( !rd2_out_last ) begin
                        state3 <= `S3_ENGINE_PROCESSING;
                    end
                end
                else begin
                    rd3_process_valid       <= 1'b0;
                end
            end
            `S3_ENGINE_PROCESSING: begin
                rd3_process_first           <= 1'b0;                    // FIRST
                rd3_process_last            <= rd3_process_next_last;   // LAST
                rd3_process_dwlen           <= rd3_process_dwlen - 1;   // LEN DEC
                rd3_process_dwaddr          <= rd3_process_dwaddr + 1;  // ADDR INC
                if ( rd3_process_next_last ) begin
                    state3 <= `S3_ENGINE_REQDATA;
                end
            end
        endcase

    assign rd2_out_rden = rd3_enable && (
        ((state3 == `S3_ENGINE_REQDATA) && (!rd2_out_valid || rd2_out_last)) ||
        ((state3 == `S3_ENGINE_PROCESSING) && rd3_process_nextnext_last));
    
    // ------------------------------------------------------------------------
    // 4: PROCESS RESPONSES:
    // ------------------------------------------------------------------------
    
    wire        rd_rsp_first    = rd_rsp_ctx[87];
    wire        rd_rsp_last     = rd_rsp_ctx[86];
    
    wire [9:0]  rd_rsp_dwlen    = rd_rsp_ctx[72:63];
    wire [11:0] rd_rsp_bc       = rd_rsp_ctx[85:74];
    wire [15:0] rd_rsp_reqid    = rd_rsp_ctx[47:32];
    wire [7:0]  rd_rsp_tag      = rd_rsp_ctx[55:48];
    wire [6:0]  rd_rsp_lowaddr  = rd_rsp_ctx[6:0];
    wire [31:0] rd_rsp_addr     = rd_rsp_ctx[31:0];
    wire [31:0] rd_rsp_data_bs  = { rd_rsp_data[7:0], rd_rsp_data[15:8], rd_rsp_data[23:16], rd_rsp_data[31:24] };
    
    // 1: 32-bit -> 128-bit state machine:
    bit [127:0] tdata;
    bit [3:0]   tkeepdw = 0;
    bit         tlast;
    bit         first   = 1;
    wire        tvalid  = tlast || tkeepdw[3];
    
    always @ ( posedge clk )
        if ( rst ) begin
            tkeepdw <= 0;
            tlast   <= 0;
            first   <= 0;
        end
        else if ( rd_rsp_valid && rd_rsp_first ) begin
            tkeepdw         <= 4'b1111;
            tlast           <= rd_rsp_last;
            first           <= 1'b1;
            tdata[31:0]     <= { 22'b0100101000000000000000, rd_rsp_dwlen };            // format, type, length
            tdata[63:32]    <= { pcie_id[7:0], pcie_id[15:8], 4'b0, rd_rsp_bc };        // pcie_id, byte_count
            tdata[95:64]    <= { rd_rsp_reqid, rd_rsp_tag, 1'b0, rd_rsp_lowaddr };      // req_id, tag, lower_addr
            tdata[127:96]   <= rd_rsp_data_bs;
        end
        else begin
            tlast   <= rd_rsp_valid && rd_rsp_last;
            tkeepdw <= tvalid ? (rd_rsp_valid ? 4'b0001 : 4'b0000) : (rd_rsp_valid ? ((tkeepdw << 1) | 1'b1) : tkeepdw);
            first   <= 0;
            if ( rd_rsp_valid ) begin
                if ( tvalid || !tkeepdw[0] )
                    tdata[31:0]   <= rd_rsp_data_bs;
                if ( !tkeepdw[1] )
                    tdata[63:32]  <= rd_rsp_data_bs;
                if ( !tkeepdw[2] )
                    tdata[95:64]  <= rd_rsp_data_bs;
                if ( !tkeepdw[3] )
                    tdata[127:96] <= rd_rsp_data_bs;   
            end
        end
    
    // 2.1 - submit to output fifo - will feed into mux/pcie core.
    fifo_134_134_clk1_bar_rdrsp i_fifo_134_134_clk1_bar_rdrsp(
        .srst           ( rst                       ),
        .clk            ( clk                       ),
        .din            ( { first, tlast, tkeepdw, tdata } ),
        .wr_en          ( tvalid                    ),
        .rd_en          ( tlps_out.tready           ),
        .dout           ( { tlps_out.tuser[0], tlps_out.tlast, tlps_out.tkeepdw, tlps_out.tdata } ),
        .full           (                           ),
        .empty          (                           ),
        .prog_empty     ( rd3_enable                ),
        .valid          ( tlps_out.tvalid           )
    );
    
    assign tlps_out.tuser[1] = tlps_out.tlast;
    assign tlps_out.tuser[8:2] = 0;
    
    // 2.2 - packet count:
    bit [10:0]  pkt_count       = 0;
    wire        pkt_count_dec   = tlps_out.tvalid && tlps_out.tlast;
    wire        pkt_count_inc   = tvalid && tlast;
    wire [10:0] pkt_count_next  = pkt_count + pkt_count_inc - pkt_count_dec;
    assign tlps_out.has_data    = (pkt_count_next > 0);
    
    always @ ( posedge clk ) begin
        pkt_count <= rst ? 0 : pkt_count_next;
    end

endmodule


// ------------------------------------------------------------------------
// Example BAR implementation that does nothing but drop any read/writes
// silently without generating a response.
// This is only recommended for placeholder designs.
// Latency = N/A.
// ------------------------------------------------------------------------
module pcileech_bar_impl_none(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    initial rd_rsp_ctx = 0;
    initial rd_rsp_data = 0;
    initial rd_rsp_valid = 0;

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of "address loopback" which can be useful
// for testing. Any read to a specific BAR address will result in the
// address as response.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_loopaddr(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input [87:0]        rd_req_ctx,
    input [31:0]        rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]      rd_req_ctx_1;
    bit [31:0]      rd_req_addr_1;
    bit             rd_req_valid_1;
    
    always @ ( posedge clk ) begin
        rd_req_ctx_1    <= rd_req_ctx;
        rd_req_addr_1   <= rd_req_addr;
        rd_req_valid_1  <= rd_req_valid;
        rd_rsp_ctx      <= rd_req_ctx_1;
        rd_rsp_data     <= rd_req_addr_1;
        rd_rsp_valid    <= rd_req_valid_1;
    end    

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of a 4kB writable initial-zero BAR.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_zerowrite4k(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]  drd_req_ctx;
    bit         drd_req_valid;
    wire [31:0] doutb;
    
    always @ ( posedge clk ) begin
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        rd_rsp_data     <= doutb; 
    end
    
    bram_bar_zero4k i_bram_bar_zero4k(
        // Port A - write:
        .addra  ( wr_addr[11:2]     ),
        .clka   ( clk               ),
        .dina   ( wr_data           ),
        .ena    ( wr_valid          ),
        .wea    ( wr_be             ),
        // Port A - read (2 CLK latency):
        .addrb  ( rd_req_addr[11:2] ),
        .clkb   ( clk               ),
        .doutb  ( doutb             ),
        .enb    ( rd_req_valid      )
    );

endmodule



// 这是一个bar2的tlp回应实现
module pcileech_bar_impl_bar2(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    input  [31:0]       base_address_register,
    // outgoing BAR read replies:
    output reg [87:0]   rd_rsp_ctx,
    output reg [31:0]   rd_rsp_data,
    output reg          rd_rsp_valid
);
                     
    reg [87:0]      drd_req_ctx;
    reg [31:0]      drd_req_addr;
    reg             drd_req_valid;
                  
    reg [31:0]      dwr_addr;
    reg [31:0]      dwr_data;
    reg             dwr_valid;
               
    reg [31:0]      data_32;
              
    time number = 0;
                  
    always @ (posedge clk) begin
        if (rst)
            number <= 0;
               
        number          <= number + 1;
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        dwr_valid       <= wr_valid;
        drd_req_addr    <= rd_req_addr;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        dwr_addr        <= wr_addr;
        dwr_data        <= wr_data;

        
        

        if (drd_req_valid) begin
            // 52104004 - 52104000 = 00000004 & FFFF = 0004
            case (({drd_req_addr[31:24], drd_req_addr[23:16], drd_req_addr[15:08], drd_req_addr[07:00]} - (base_address_register & 32'hFFFFFFF0)) & 32'h0FFF)
                16'h0000 : rd_rsp_data <= 32'h03B4BE60;
                16'h0004 : rd_rsp_data <= 32'h00006EF0;
                16'h0008 : rd_rsp_data <= 32'h80000040;
                16'h000C : rd_rsp_data <= 32'h00000080;
                16'h0010 : rd_rsp_data <= 32'h9A086C00;
                16'h0014 : rd_rsp_data <= 32'h00000001;
                16'h0018 : rd_rsp_data <= 32'h00460807;
                16'h0020 : rd_rsp_data <= 32'h9A087000;
                16'h0024 : rd_rsp_data <= 32'h00000001;
                16'h0028 : rd_rsp_data <= 32'h9A0BD000;
                16'h002C : rd_rsp_data <= 32'h00000001;
                16'h003C : rd_rsp_data <= 32'h00210021;
                16'h0040 : rd_rsp_data <= 32'h54100800;
                16'h0044 : rd_rsp_data <= 32'h01020F00;
                16'h0050 : rd_rsp_data <= 32'hBCCF0010;
                16'h0054 : rd_rsp_data <= 32'h01031160;
                16'h0064 : rd_rsp_data <= 32'h27FFFF01;
                16'h0068 : rd_rsp_data <= 32'h0000870C;
                16'h006C : rd_rsp_data <= 32'hF0C00004;
                16'h0070 : rd_rsp_data <= 32'h00000001;
                16'h0074 : rd_rsp_data <= 32'h0000F2FC;
                16'h0078 : rd_rsp_data <= 32'h00000007;
                16'h0080 : rd_rsp_data <= 32'h0001068B;
                16'h00B4 : rd_rsp_data <= 32'h00010000;
                16'h00B8 : rd_rsp_data <= 32'hD2017989;
                16'h00D0 : rd_rsp_data <= 32'h320000E1;
                16'h00D4 : rd_rsp_data <= 32'h0000000E;
                16'h00D8 : rd_rsp_data <= 32'h05F30000;
                16'h00DC : rd_rsp_data <= 32'h007DCC83;
                16'h00E0 : rd_rsp_data <= 32'h00002060;
                16'h00E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h00E8 : rd_rsp_data <= 32'h00000001;
                16'h00EC : rd_rsp_data <= 32'h0000003F;
                16'h00F0 : rd_rsp_data <= 32'h0048803F;
                16'h00F8 : rd_rsp_data <= 32'h00000003;
                16'h0100 : rd_rsp_data <= 32'h03B4BE60;
                16'h0104 : rd_rsp_data <= 32'h00006EF0;
                16'h0108 : rd_rsp_data <= 32'h80000040;
                16'h010C : rd_rsp_data <= 32'h00000080;
                16'h0110 : rd_rsp_data <= 32'h9A086C00;
                16'h0114 : rd_rsp_data <= 32'h00000001;
                16'h0118 : rd_rsp_data <= 32'h00460807;
                16'h0120 : rd_rsp_data <= 32'h9A087000;
                16'h0124 : rd_rsp_data <= 32'h00000001;
                16'h0128 : rd_rsp_data <= 32'h9A0BD000;
                16'h012C : rd_rsp_data <= 32'h00000001;
                16'h0140 : rd_rsp_data <= 32'h54100800;
                16'h0144 : rd_rsp_data <= 32'h01020F00;
                16'h0150 : rd_rsp_data <= 32'hBCCF0010;
                16'h0154 : rd_rsp_data <= 32'h01031160;
                16'h0164 : rd_rsp_data <= 32'h27FFFF01;
                16'h0168 : rd_rsp_data <= 32'h0000870C;
                16'h016C : rd_rsp_data <= 32'hF0C00004;
                16'h0170 : rd_rsp_data <= 32'h00000001;
                16'h0174 : rd_rsp_data <= 32'h0000F2FC;
                16'h0178 : rd_rsp_data <= 32'h00000007;
                16'h0180 : rd_rsp_data <= 32'h0001068B;
                16'h01B4 : rd_rsp_data <= 32'h00010000;
                16'h01B8 : rd_rsp_data <= 32'hD2017989;
                16'h01D0 : rd_rsp_data <= 32'h320000E1;
                16'h01D4 : rd_rsp_data <= 32'h0000000E;
                16'h01D8 : rd_rsp_data <= 32'h05F30000;
                16'h01DC : rd_rsp_data <= 32'h007DCC83;
                16'h01E0 : rd_rsp_data <= 32'h00002060;
                16'h01E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h01E8 : rd_rsp_data <= 32'h00000001;
                16'h01EC : rd_rsp_data <= 32'h0000003F;
                16'h01F0 : rd_rsp_data <= 32'h0048803F;
                16'h01F8 : rd_rsp_data <= 32'h00000003;
                16'h0200 : rd_rsp_data <= 32'h03B4BE60;
                16'h0204 : rd_rsp_data <= 32'h00006EF0;
                16'h0208 : rd_rsp_data <= 32'h80000040;
                16'h020C : rd_rsp_data <= 32'h00000080;
                16'h0210 : rd_rsp_data <= 32'h9A086C00;
                16'h0214 : rd_rsp_data <= 32'h00000001;
                16'h0218 : rd_rsp_data <= 32'h00460807;
                16'h0220 : rd_rsp_data <= 32'h9A087000;
                16'h0224 : rd_rsp_data <= 32'h00000001;
                16'h0228 : rd_rsp_data <= 32'h9A0BD000;
                16'h022C : rd_rsp_data <= 32'h00000001;
                16'h0240 : rd_rsp_data <= 32'h54100800;
                16'h0244 : rd_rsp_data <= 32'h01020F00;
                16'h0250 : rd_rsp_data <= 32'hBCCF0010;
                16'h0254 : rd_rsp_data <= 32'h01031160;
                16'h0264 : rd_rsp_data <= 32'h27FFFF01;
                16'h0268 : rd_rsp_data <= 32'h0000870C;
                16'h026C : rd_rsp_data <= 32'hF0C00004;
                16'h0270 : rd_rsp_data <= 32'h00000001;
                16'h0274 : rd_rsp_data <= 32'h0000F2FC;
                16'h0278 : rd_rsp_data <= 32'h00000007;
                16'h0280 : rd_rsp_data <= 32'h0001068B;
                16'h02B4 : rd_rsp_data <= 32'h00010000;
                16'h02B8 : rd_rsp_data <= 32'hD2017989;
                16'h02D0 : rd_rsp_data <= 32'h320000E1;
                16'h02D4 : rd_rsp_data <= 32'h0000000E;
                16'h02D8 : rd_rsp_data <= 32'h05F30000;
                16'h02DC : rd_rsp_data <= 32'h007DCC83;
                16'h02E0 : rd_rsp_data <= 32'h00002060;
                16'h02E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h02E8 : rd_rsp_data <= 32'h00000001;
                16'h02EC : rd_rsp_data <= 32'h0000003F;
                16'h02F0 : rd_rsp_data <= 32'h0048803F;
                16'h02F8 : rd_rsp_data <= 32'h00000003;
                16'h0300 : rd_rsp_data <= 32'h03B4BE60;
                16'h0304 : rd_rsp_data <= 32'h00006EF0;
                16'h0308 : rd_rsp_data <= 32'h80000040;
                16'h030C : rd_rsp_data <= 32'h00000080;
                16'h0310 : rd_rsp_data <= 32'h9A086C00;
                16'h0314 : rd_rsp_data <= 32'h00000001;
                16'h0318 : rd_rsp_data <= 32'h00460807;
                16'h0320 : rd_rsp_data <= 32'h9A087000;
                16'h0324 : rd_rsp_data <= 32'h00000001;
                16'h0328 : rd_rsp_data <= 32'h9A0BD000;
                16'h032C : rd_rsp_data <= 32'h00000001;
                16'h0340 : rd_rsp_data <= 32'h54100800;
                16'h0344 : rd_rsp_data <= 32'h01020F00;
                16'h0350 : rd_rsp_data <= 32'hBCCF0010;
                16'h0354 : rd_rsp_data <= 32'h01031160;
                16'h0364 : rd_rsp_data <= 32'h27FFFF01;
                16'h0368 : rd_rsp_data <= 32'h0000870C;
                16'h036C : rd_rsp_data <= 32'hF0C00004;
                16'h0370 : rd_rsp_data <= 32'h00000001;
                16'h0374 : rd_rsp_data <= 32'h0000F2FC;
                16'h0378 : rd_rsp_data <= 32'h00000007;
                16'h0380 : rd_rsp_data <= 32'h0001068B;
                16'h03B4 : rd_rsp_data <= 32'h00010000;
                16'h03B8 : rd_rsp_data <= 32'hD2017989;
                16'h03D0 : rd_rsp_data <= 32'h320000E1;
                16'h03D4 : rd_rsp_data <= 32'h0000000E;
                16'h03D8 : rd_rsp_data <= 32'h05F30000;
                16'h03DC : rd_rsp_data <= 32'h007DCC83;
                16'h03E0 : rd_rsp_data <= 32'h00002060;
                16'h03E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h03E8 : rd_rsp_data <= 32'h00000001;
                16'h03EC : rd_rsp_data <= 32'h0000003F;
                16'h03F0 : rd_rsp_data <= 32'h0048803F;
                16'h03F8 : rd_rsp_data <= 32'h00000003;
                16'h0400 : rd_rsp_data <= 32'h03B4BE60;
                16'h0404 : rd_rsp_data <= 32'h00006EF0;
                16'h0408 : rd_rsp_data <= 32'h80000040;
                16'h040C : rd_rsp_data <= 32'h00000080;
                16'h0410 : rd_rsp_data <= 32'h9A086C00;
                16'h0414 : rd_rsp_data <= 32'h00000001;
                16'h0418 : rd_rsp_data <= 32'h00460807;
                16'h0420 : rd_rsp_data <= 32'h9A087000;
                16'h0424 : rd_rsp_data <= 32'h00000001;
                16'h0428 : rd_rsp_data <= 32'h9A0BD000;
                16'h042C : rd_rsp_data <= 32'h00000001;
                16'h0440 : rd_rsp_data <= 32'h54100800;
                16'h0444 : rd_rsp_data <= 32'h01020F00;
                16'h0450 : rd_rsp_data <= 32'hBCCF0010;
                16'h0454 : rd_rsp_data <= 32'h01031160;
                16'h0464 : rd_rsp_data <= 32'h27FFFF01;
                16'h0468 : rd_rsp_data <= 32'h0000870C;
                16'h046C : rd_rsp_data <= 32'hF0C00004;
                16'h0470 : rd_rsp_data <= 32'h00000001;
                16'h0474 : rd_rsp_data <= 32'h0000F2FC;
                16'h0478 : rd_rsp_data <= 32'h00000007;
                16'h0480 : rd_rsp_data <= 32'h0001068B;
                16'h04B4 : rd_rsp_data <= 32'h00010000;
                16'h04B8 : rd_rsp_data <= 32'hD2017989;
                16'h04D0 : rd_rsp_data <= 32'h320000E1;
                16'h04D4 : rd_rsp_data <= 32'h0000000E;
                16'h04D8 : rd_rsp_data <= 32'h05F30000;
                16'h04DC : rd_rsp_data <= 32'h007DCC83;
                16'h04E0 : rd_rsp_data <= 32'h00002060;
                16'h04E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h04E8 : rd_rsp_data <= 32'h00000001;
                16'h04EC : rd_rsp_data <= 32'h0000003F;
                16'h04F0 : rd_rsp_data <= 32'h0048803F;
                16'h04F8 : rd_rsp_data <= 32'h00000003;
                16'h0500 : rd_rsp_data <= 32'h03B4BE60;
                16'h0504 : rd_rsp_data <= 32'h00006EF0;
                16'h0508 : rd_rsp_data <= 32'h80000040;
                16'h050C : rd_rsp_data <= 32'h00000080;
                16'h0510 : rd_rsp_data <= 32'h9A086C00;
                16'h0514 : rd_rsp_data <= 32'h00000001;
                16'h0518 : rd_rsp_data <= 32'h00460807;
                16'h0520 : rd_rsp_data <= 32'h9A087000;
                16'h0524 : rd_rsp_data <= 32'h00000001;
                16'h0528 : rd_rsp_data <= 32'h9A0BD000;
                16'h052C : rd_rsp_data <= 32'h00000001;
                16'h0540 : rd_rsp_data <= 32'h54100800;
                16'h0544 : rd_rsp_data <= 32'h01020F00;
                16'h0550 : rd_rsp_data <= 32'hBCCF0010;
                16'h0554 : rd_rsp_data <= 32'h01031160;
                16'h0564 : rd_rsp_data <= 32'h27FFFF01;
                16'h0568 : rd_rsp_data <= 32'h0000870C;
                16'h056C : rd_rsp_data <= 32'hF0C00004;
                16'h0570 : rd_rsp_data <= 32'h00000001;
                16'h0574 : rd_rsp_data <= 32'h0000F2FC;
                16'h0578 : rd_rsp_data <= 32'h00000007;
                16'h0580 : rd_rsp_data <= 32'h0001068B;
                16'h05B4 : rd_rsp_data <= 32'h00010000;
                16'h05B8 : rd_rsp_data <= 32'hD2017989;
                16'h05D0 : rd_rsp_data <= 32'h320000E1;
                16'h05D4 : rd_rsp_data <= 32'h0000000E;
                16'h05D8 : rd_rsp_data <= 32'h05F30000;
                16'h05DC : rd_rsp_data <= 32'h007DCC83;
                16'h05E0 : rd_rsp_data <= 32'h00002060;
                16'h05E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h05E8 : rd_rsp_data <= 32'h00000001;
                16'h05EC : rd_rsp_data <= 32'h0000003F;
                16'h05F0 : rd_rsp_data <= 32'h0048803F;
                16'h05F8 : rd_rsp_data <= 32'h00000003;
                16'h0600 : rd_rsp_data <= 32'h03B4BE60;
                16'h0604 : rd_rsp_data <= 32'h00006EF0;
                16'h0608 : rd_rsp_data <= 32'h80000040;
                16'h060C : rd_rsp_data <= 32'h00000080;
                16'h0610 : rd_rsp_data <= 32'h9A086C00;
                16'h0614 : rd_rsp_data <= 32'h00000001;
                16'h0618 : rd_rsp_data <= 32'h00460807;
                16'h0620 : rd_rsp_data <= 32'h9A087000;
                16'h0624 : rd_rsp_data <= 32'h00000001;
                16'h0628 : rd_rsp_data <= 32'h9A0BD000;
                16'h062C : rd_rsp_data <= 32'h00000001;
                16'h0640 : rd_rsp_data <= 32'h54100800;
                16'h0644 : rd_rsp_data <= 32'h01020F00;
                16'h0650 : rd_rsp_data <= 32'hBCCF0010;
                16'h0654 : rd_rsp_data <= 32'h01031160;
                16'h0664 : rd_rsp_data <= 32'h27FFFF01;
                16'h0668 : rd_rsp_data <= 32'h0000870C;
                16'h066C : rd_rsp_data <= 32'hF0C00004;
                16'h0670 : rd_rsp_data <= 32'h00000001;
                16'h0674 : rd_rsp_data <= 32'h0000F2FC;
                16'h0678 : rd_rsp_data <= 32'h00000007;
                16'h0680 : rd_rsp_data <= 32'h0001068B;
                16'h06B4 : rd_rsp_data <= 32'h00010000;
                16'h06B8 : rd_rsp_data <= 32'hD2017989;
                16'h06D0 : rd_rsp_data <= 32'h320000E1;
                16'h06D4 : rd_rsp_data <= 32'h0000000E;
                16'h06D8 : rd_rsp_data <= 32'h05F30000;
                16'h06DC : rd_rsp_data <= 32'h007DCC83;
                16'h06E0 : rd_rsp_data <= 32'h00002060;
                16'h06E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h06E8 : rd_rsp_data <= 32'h00000001;
                16'h06EC : rd_rsp_data <= 32'h0000003F;
                16'h06F0 : rd_rsp_data <= 32'h0048803F;
                16'h06F8 : rd_rsp_data <= 32'h00000003;
                16'h0700 : rd_rsp_data <= 32'h03B4BE60;
                16'h0704 : rd_rsp_data <= 32'h00006EF0;
                16'h0708 : rd_rsp_data <= 32'h80000040;
                16'h070C : rd_rsp_data <= 32'h00000080;
                16'h0710 : rd_rsp_data <= 32'h9A086C00;
                16'h0714 : rd_rsp_data <= 32'h00000001;
                16'h0718 : rd_rsp_data <= 32'h00460807;
                16'h0720 : rd_rsp_data <= 32'h9A087000;
                16'h0724 : rd_rsp_data <= 32'h00000001;
                16'h0728 : rd_rsp_data <= 32'h9A0BD000;
                16'h072C : rd_rsp_data <= 32'h00000001;
                16'h0740 : rd_rsp_data <= 32'h54100800;
                16'h0744 : rd_rsp_data <= 32'h01020F00;
                16'h0750 : rd_rsp_data <= 32'hBCCF0010;
                16'h0754 : rd_rsp_data <= 32'h01031160;
                16'h0764 : rd_rsp_data <= 32'h27FFFF01;
                16'h0768 : rd_rsp_data <= 32'h0000870C;
                16'h076C : rd_rsp_data <= 32'hF0C00004;
                16'h0770 : rd_rsp_data <= 32'h00000001;
                16'h0774 : rd_rsp_data <= 32'h0000F2FC;
                16'h0778 : rd_rsp_data <= 32'h00000007;
                16'h0780 : rd_rsp_data <= 32'h0001068B;
                16'h07B4 : rd_rsp_data <= 32'h00010000;
                16'h07B8 : rd_rsp_data <= 32'hD2017989;
                16'h07D0 : rd_rsp_data <= 32'h320000E1;
                16'h07D4 : rd_rsp_data <= 32'h0000000E;
                16'h07D8 : rd_rsp_data <= 32'h05F30000;
                16'h07DC : rd_rsp_data <= 32'h007DCC83;
                16'h07E0 : rd_rsp_data <= 32'h00002060;
                16'h07E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h07E8 : rd_rsp_data <= 32'h00000001;
                16'h07EC : rd_rsp_data <= 32'h0000003F;
                16'h07F0 : rd_rsp_data <= 32'h0048803F;
                16'h07F8 : rd_rsp_data <= 32'h00000003;
                16'h0800 : rd_rsp_data <= 32'h03B4BE60;
                16'h0804 : rd_rsp_data <= 32'h00006EF0;
                16'h0808 : rd_rsp_data <= 32'h80000040;
                16'h080C : rd_rsp_data <= 32'h00000080;
                16'h0810 : rd_rsp_data <= 32'h9A086C00;
                16'h0814 : rd_rsp_data <= 32'h00000001;
                16'h0818 : rd_rsp_data <= 32'h00460807;
                16'h0820 : rd_rsp_data <= 32'h9A087000;
                16'h0824 : rd_rsp_data <= 32'h00000001;
                16'h0828 : rd_rsp_data <= 32'h9A0BD000;
                16'h082C : rd_rsp_data <= 32'h00000001;
                16'h0840 : rd_rsp_data <= 32'h54100800;
                16'h0844 : rd_rsp_data <= 32'h01020F00;
                16'h0850 : rd_rsp_data <= 32'hBCCF0010;
                16'h0854 : rd_rsp_data <= 32'h01031160;
                16'h0864 : rd_rsp_data <= 32'h27FFFF01;
                16'h0868 : rd_rsp_data <= 32'h0000870C;
                16'h086C : rd_rsp_data <= 32'hF0C00004;
                16'h0870 : rd_rsp_data <= 32'h00000001;
                16'h0874 : rd_rsp_data <= 32'h0000F2FC;
                16'h0878 : rd_rsp_data <= 32'h00000007;
                16'h0880 : rd_rsp_data <= 32'h0001068B;
                16'h08B4 : rd_rsp_data <= 32'h00010000;
                16'h08B8 : rd_rsp_data <= 32'hD2017989;
                16'h08D0 : rd_rsp_data <= 32'h320000E1;
                16'h08D4 : rd_rsp_data <= 32'h0000000E;
                16'h08D8 : rd_rsp_data <= 32'h05F30000;
                16'h08DC : rd_rsp_data <= 32'h007DCC83;
                16'h08E0 : rd_rsp_data <= 32'h00002060;
                16'h08E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h08E8 : rd_rsp_data <= 32'h00000001;
                16'h08EC : rd_rsp_data <= 32'h0000003F;
                16'h08F0 : rd_rsp_data <= 32'h0048803F;
                16'h08F8 : rd_rsp_data <= 32'h00000003;
                16'h0900 : rd_rsp_data <= 32'h03B4BE60;
                16'h0904 : rd_rsp_data <= 32'h00006EF0;
                16'h0908 : rd_rsp_data <= 32'h80000040;
                16'h090C : rd_rsp_data <= 32'h00000080;
                16'h0910 : rd_rsp_data <= 32'h9A086C00;
                16'h0914 : rd_rsp_data <= 32'h00000001;
                16'h0918 : rd_rsp_data <= 32'h00460807;
                16'h0920 : rd_rsp_data <= 32'h9A087000;
                16'h0924 : rd_rsp_data <= 32'h00000001;
                16'h0928 : rd_rsp_data <= 32'h9A0BD000;
                16'h092C : rd_rsp_data <= 32'h00000001;
                16'h0940 : rd_rsp_data <= 32'h54100800;
                16'h0944 : rd_rsp_data <= 32'h01020F00;
                16'h0950 : rd_rsp_data <= 32'hBCCF0010;
                16'h0954 : rd_rsp_data <= 32'h01031160;
                16'h0964 : rd_rsp_data <= 32'h27FFFF01;
                16'h0968 : rd_rsp_data <= 32'h0000870C;
                16'h096C : rd_rsp_data <= 32'hF0C00004;
                16'h0970 : rd_rsp_data <= 32'h00000001;
                16'h0974 : rd_rsp_data <= 32'h0000F2FC;
                16'h0978 : rd_rsp_data <= 32'h00000007;
                16'h0980 : rd_rsp_data <= 32'h0001068B;
                16'h09B4 : rd_rsp_data <= 32'h00010000;
                16'h09B8 : rd_rsp_data <= 32'hD2017989;
                16'h09D0 : rd_rsp_data <= 32'h320000E1;
                16'h09D4 : rd_rsp_data <= 32'h0000000E;
                16'h09D8 : rd_rsp_data <= 32'h05F30000;
                16'h09DC : rd_rsp_data <= 32'h007DCC83;
                16'h09E0 : rd_rsp_data <= 32'h00002060;
                16'h09E4 : rd_rsp_data <= 32'h9A0C0000;
                16'h09E8 : rd_rsp_data <= 32'h00000001;
                16'h09EC : rd_rsp_data <= 32'h0000003F;
                16'h09F0 : rd_rsp_data <= 32'h0048803F;
                16'h09F8 : rd_rsp_data <= 32'h00000003;
                16'h0A00 : rd_rsp_data <= 32'h03B4BE60;
                16'h0A04 : rd_rsp_data <= 32'h00006EF0;
                16'h0A08 : rd_rsp_data <= 32'h80000040;
                16'h0A0C : rd_rsp_data <= 32'h00000080;
                16'h0A10 : rd_rsp_data <= 32'h9A086C00;
                16'h0A14 : rd_rsp_data <= 32'h00000001;
                16'h0A18 : rd_rsp_data <= 32'h00460807;
                16'h0A20 : rd_rsp_data <= 32'h9A087000;
                16'h0A24 : rd_rsp_data <= 32'h00000001;
                16'h0A28 : rd_rsp_data <= 32'h9A0BD000;
                16'h0A2C : rd_rsp_data <= 32'h00000001;
                16'h0A40 : rd_rsp_data <= 32'h54100800;
                16'h0A44 : rd_rsp_data <= 32'h01020F00;
                16'h0A50 : rd_rsp_data <= 32'hBCCF0010;
                16'h0A54 : rd_rsp_data <= 32'h01031160;
                16'h0A64 : rd_rsp_data <= 32'h27FFFF01;
                16'h0A68 : rd_rsp_data <= 32'h0000870C;
                16'h0A6C : rd_rsp_data <= 32'hF0C00004;
                16'h0A70 : rd_rsp_data <= 32'h00000001;
                16'h0A74 : rd_rsp_data <= 32'h0000F2FC;
                16'h0A78 : rd_rsp_data <= 32'h00000007;
                16'h0A80 : rd_rsp_data <= 32'h0001068B;
                16'h0AB4 : rd_rsp_data <= 32'h00010000;
                16'h0AB8 : rd_rsp_data <= 32'hD2017989;
                16'h0AD0 : rd_rsp_data <= 32'h320000E1;
                16'h0AD4 : rd_rsp_data <= 32'h0000000E;
                16'h0AD8 : rd_rsp_data <= 32'h05F30000;
                16'h0ADC : rd_rsp_data <= 32'h007DCC83;
                16'h0AE0 : rd_rsp_data <= 32'h00002060;
                16'h0AE4 : rd_rsp_data <= 32'h9A0C0000;
                16'h0AE8 : rd_rsp_data <= 32'h00000001;
                16'h0AEC : rd_rsp_data <= 32'h0000003F;
                16'h0AF0 : rd_rsp_data <= 32'h0048803F;
                16'h0AF8 : rd_rsp_data <= 32'h00000003;
                16'h0B00 : rd_rsp_data <= 32'h03B4BE60;
                16'h0B04 : rd_rsp_data <= 32'h00006EF0;
                16'h0B08 : rd_rsp_data <= 32'h80000040;
                16'h0B0C : rd_rsp_data <= 32'h00000080;
                16'h0B10 : rd_rsp_data <= 32'h9A086C00;
                16'h0B14 : rd_rsp_data <= 32'h00000001;
                16'h0B18 : rd_rsp_data <= 32'h00460807;
                16'h0B20 : rd_rsp_data <= 32'h9A087000;
                16'h0B24 : rd_rsp_data <= 32'h00000001;
                16'h0B28 : rd_rsp_data <= 32'h9A0BD000;
                16'h0B2C : rd_rsp_data <= 32'h00000001;
                16'h0B40 : rd_rsp_data <= 32'h54100800;
                16'h0B44 : rd_rsp_data <= 32'h01020F00;
                16'h0B50 : rd_rsp_data <= 32'hBCCF0010;
                16'h0B54 : rd_rsp_data <= 32'h01031160;
                16'h0B64 : rd_rsp_data <= 32'h27FFFF01;
                16'h0B68 : rd_rsp_data <= 32'h0000870C;
                16'h0B6C : rd_rsp_data <= 32'hF0C00004;
                16'h0B70 : rd_rsp_data <= 32'h00000001;
                16'h0B74 : rd_rsp_data <= 32'h0000F2FC;
                16'h0B78 : rd_rsp_data <= 32'h00000007;
                16'h0B80 : rd_rsp_data <= 32'h0001068B;
                16'h0BB4 : rd_rsp_data <= 32'h00010000;
                16'h0BB8 : rd_rsp_data <= 32'hD2017989;
                16'h0BD0 : rd_rsp_data <= 32'h320000E1;
                16'h0BD4 : rd_rsp_data <= 32'h0000000E;
                16'h0BD8 : rd_rsp_data <= 32'h05F30000;
                16'h0BDC : rd_rsp_data <= 32'h007DCC83;
                16'h0BE0 : rd_rsp_data <= 32'h00002060;
                16'h0BE4 : rd_rsp_data <= 32'h9A0C0000;
                16'h0BE8 : rd_rsp_data <= 32'h00000001;
                16'h0BEC : rd_rsp_data <= 32'h0000003F;
                16'h0BF0 : rd_rsp_data <= 32'h0048803F;
                16'h0BF8 : rd_rsp_data <= 32'h00000003;
                16'h0C00 : rd_rsp_data <= 32'h03B4BE60;
                16'h0C04 : rd_rsp_data <= 32'h00006EF0;
                16'h0C08 : rd_rsp_data <= 32'h80000040;
                16'h0C0C : rd_rsp_data <= 32'h00000080;
                16'h0C10 : rd_rsp_data <= 32'h9A086C00;
                16'h0C14 : rd_rsp_data <= 32'h00000001;
                16'h0C18 : rd_rsp_data <= 32'h00460807;
                16'h0C20 : rd_rsp_data <= 32'h9A087000;
                16'h0C24 : rd_rsp_data <= 32'h00000001;
                16'h0C28 : rd_rsp_data <= 32'h9A0BD000;
                16'h0C2C : rd_rsp_data <= 32'h00000001;
                16'h0C40 : rd_rsp_data <= 32'h54100800;
                16'h0C44 : rd_rsp_data <= 32'h01020F00;
                16'h0C50 : rd_rsp_data <= 32'hBCCF0010;
                16'h0C54 : rd_rsp_data <= 32'h01031160;
                16'h0C64 : rd_rsp_data <= 32'h27FFFF01;
                16'h0C68 : rd_rsp_data <= 32'h0000870C;
                16'h0C6C : rd_rsp_data <= 32'hF0C00004;
                16'h0C70 : rd_rsp_data <= 32'h00000001;
                16'h0C74 : rd_rsp_data <= 32'h0000F2FC;
                16'h0C78 : rd_rsp_data <= 32'h00000007;
                16'h0C80 : rd_rsp_data <= 32'h0001068B;
                16'h0CB4 : rd_rsp_data <= 32'h00010000;
                16'h0CB8 : rd_rsp_data <= 32'hD2017989;
                16'h0CD0 : rd_rsp_data <= 32'h320000E1;
                16'h0CD4 : rd_rsp_data <= 32'h0000000E;
                16'h0CD8 : rd_rsp_data <= 32'h05F30000;
                16'h0CDC : rd_rsp_data <= 32'h007DCC83;
                16'h0CE0 : rd_rsp_data <= 32'h00002060;
                16'h0CE4 : rd_rsp_data <= 32'h9A0C0000;
                16'h0CE8 : rd_rsp_data <= 32'h00000001;
                16'h0CEC : rd_rsp_data <= 32'h0000003F;
                16'h0CF0 : rd_rsp_data <= 32'h0048803F;
                16'h0CF8 : rd_rsp_data <= 32'h00000003;
                16'h0D00 : rd_rsp_data <= 32'h03B4BE60;
                16'h0D04 : rd_rsp_data <= 32'h00006EF0;
                16'h0D08 : rd_rsp_data <= 32'h80000040;
                16'h0D0C : rd_rsp_data <= 32'h00000080;
                16'h0D10 : rd_rsp_data <= 32'h9A086C00;
                16'h0D14 : rd_rsp_data <= 32'h00000001;
                16'h0D18 : rd_rsp_data <= 32'h00460807;
                16'h0D20 : rd_rsp_data <= 32'h9A087000;
                16'h0D24 : rd_rsp_data <= 32'h00000001;
                16'h0D28 : rd_rsp_data <= 32'h9A0BD000;
                16'h0D2C : rd_rsp_data <= 32'h00000001;
                16'h0D40 : rd_rsp_data <= 32'h54100800;
                16'h0D44 : rd_rsp_data <= 32'h01020F00;
                16'h0D50 : rd_rsp_data <= 32'hBCCF0010;
                16'h0D54 : rd_rsp_data <= 32'h01031160;
                16'h0D64 : rd_rsp_data <= 32'h27FFFF01;
                16'h0D68 : rd_rsp_data <= 32'h0000870C;
                16'h0D6C : rd_rsp_data <= 32'hF0C00004;
                16'h0D70 : rd_rsp_data <= 32'h00000001;
                16'h0D74 : rd_rsp_data <= 32'h0000F2FC;
                16'h0D78 : rd_rsp_data <= 32'h00000007;
                16'h0D80 : rd_rsp_data <= 32'h0001068B;
                16'h0DB4 : rd_rsp_data <= 32'h00010000;
                16'h0DB8 : rd_rsp_data <= 32'hD2017989;
                16'h0DD0 : rd_rsp_data <= 32'h320000E1;
                16'h0DD4 : rd_rsp_data <= 32'h0000000E;
                16'h0DD8 : rd_rsp_data <= 32'h05F30000;
                16'h0DDC : rd_rsp_data <= 32'h007DCC83;
                16'h0DE0 : rd_rsp_data <= 32'h00002060;
                16'h0DE4 : rd_rsp_data <= 32'h9A0C0000;
                16'h0DE8 : rd_rsp_data <= 32'h00000001;
                16'h0DEC : rd_rsp_data <= 32'h0000003F;
                16'h0DF0 : rd_rsp_data <= 32'h0048803F;
                16'h0DF8 : rd_rsp_data <= 32'h00000003;
                16'h0E00 : rd_rsp_data <= 32'h03B4BE60;
                16'h0E04 : rd_rsp_data <= 32'h00006EF0;
                16'h0E08 : rd_rsp_data <= 32'h80000040;
                16'h0E0C : rd_rsp_data <= 32'h00000080;
                16'h0E10 : rd_rsp_data <= 32'h9A086C00;
                16'h0E14 : rd_rsp_data <= 32'h00000001;
                16'h0E18 : rd_rsp_data <= 32'h00460807;
                16'h0E20 : rd_rsp_data <= 32'h9A087000;
                16'h0E24 : rd_rsp_data <= 32'h00000001;
                16'h0E28 : rd_rsp_data <= 32'h9A0BD000;
                16'h0E2C : rd_rsp_data <= 32'h00000001;
                16'h0E40 : rd_rsp_data <= 32'h54100800;
                16'h0E44 : rd_rsp_data <= 32'h01020F00;
                16'h0E50 : rd_rsp_data <= 32'hBCCF0010;
                16'h0E54 : rd_rsp_data <= 32'h01031160;
                16'h0E64 : rd_rsp_data <= 32'h27FFFF01;
                16'h0E68 : rd_rsp_data <= 32'h0000870C;
                16'h0E6C : rd_rsp_data <= 32'hF0C00004;
                16'h0E70 : rd_rsp_data <= 32'h00000001;
                16'h0E74 : rd_rsp_data <= 32'h0000F2FC;
                16'h0E78 : rd_rsp_data <= 32'h00000007;
                16'h0E80 : rd_rsp_data <= 32'h0001068B;
                16'h0EB4 : rd_rsp_data <= 32'h00010000;
                16'h0EB8 : rd_rsp_data <= 32'hD2017989;
                16'h0ED0 : rd_rsp_data <= 32'h320000E1;
                16'h0ED4 : rd_rsp_data <= 32'h0000000E;
                16'h0ED8 : rd_rsp_data <= 32'h05F30000;
                16'h0EDC : rd_rsp_data <= 32'h007DCC83;
                16'h0EE0 : rd_rsp_data <= 32'h00002060;
                16'h0EE4 : rd_rsp_data <= 32'h9A0C0000;
                16'h0EE8 : rd_rsp_data <= 32'h00000001;
                16'h0EEC : rd_rsp_data <= 32'h0000003F;
                16'h0EF0 : rd_rsp_data <= 32'h0048803F;
                16'h0EF8 : rd_rsp_data <= 32'h00000003;
                16'h0F00 : rd_rsp_data <= 32'h03B4BE60;
                16'h0F04 : rd_rsp_data <= 32'h00006EF0;
                16'h0F08 : rd_rsp_data <= 32'h80000040;
                16'h0F0C : rd_rsp_data <= 32'h00000080;
                16'h0F10 : rd_rsp_data <= 32'h9A086C00;
                16'h0F14 : rd_rsp_data <= 32'h00000001;
                16'h0F18 : rd_rsp_data <= 32'h00460807;
                16'h0F20 : rd_rsp_data <= 32'h9A087000;
                16'h0F24 : rd_rsp_data <= 32'h00000001;
                16'h0F28 : rd_rsp_data <= 32'h9A0BD000;
                16'h0F2C : rd_rsp_data <= 32'h00000001;
                16'h0F40 : rd_rsp_data <= 32'h54100800;
                16'h0F44 : rd_rsp_data <= 32'h01020F00;
                16'h0F50 : rd_rsp_data <= 32'hBCCF0010;
                16'h0F54 : rd_rsp_data <= 32'h01031160;
                16'h0F64 : rd_rsp_data <= 32'h27FFFF01;
                16'h0F68 : rd_rsp_data <= 32'h0000870C;
                16'h0F6C : rd_rsp_data <= 32'hF0C00004;
                16'h0F70 : rd_rsp_data <= 32'h00000001;
                16'h0F74 : rd_rsp_data <= 32'h0000F2FC;
                16'h0F78 : rd_rsp_data <= 32'h00000007;
                16'h0F80 : rd_rsp_data <= 32'h0001068B;
                16'h0FB4 : rd_rsp_data <= 32'h00010000;
                16'h0FB8 : rd_rsp_data <= 32'hD2017989;
                16'h0FD0 : rd_rsp_data <= 32'h320000E1;
                16'h0FD4 : rd_rsp_data <= 32'h0000000E;
                16'h0FD8 : rd_rsp_data <= 32'h05F30000;
                16'h0FDC : rd_rsp_data <= 32'h007DCC83;
                16'h0FE0 : rd_rsp_data <= 32'h00002060;
                16'h0FE4 : rd_rsp_data <= 32'h9A0C0000;
                16'h0FE8 : rd_rsp_data <= 32'h00000001;
                16'h0FEC : rd_rsp_data <= 32'h0000003F;
                16'h0FF0 : rd_rsp_data <= 32'h0048803F;
                16'h0FF8 : rd_rsp_data <= 32'h00000003;
                default: rd_rsp_data <= 32'h00000000;
            endcase
        end else if (dwr_valid) begin
            case (({dwr_addr[31:24], dwr_addr[23:16], dwr_addr[15:08], dwr_addr[07:00]} - (base_address_register & 32'hFFFFFFF0)) & 32'hFFFF)
                //Dont be scared
            endcase
        end else begin
            rd_rsp_data <= 32'h00000000;
        end
    end
            
endmodule



// 这是bar4的tlp回应实现
module pcileech_bar_impl_bar4(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    input  [31:0]       base_address_register,
    // outgoing BAR read replies:
    output reg [87:0]   rd_rsp_ctx,
    output reg [31:0]   rd_rsp_data,
    output reg          rd_rsp_valid
);
                     
    reg [87:0]      drd_req_ctx;
    reg [31:0]      drd_req_addr;
    reg             drd_req_valid;
                  
    reg [31:0]      dwr_addr;
    reg [31:0]      dwr_data;
    reg             dwr_valid;
               
    reg [31:0]      data_32;
              
    time number = 0;
                  
    always @ (posedge clk) begin
        if (rst)
            number <= 0;
               
        number          <= number + 1;
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        dwr_valid       <= wr_valid;
        drd_req_addr    <= rd_req_addr;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        dwr_addr        <= wr_addr;
        dwr_data        <= wr_data;

        if (drd_req_valid) begin
            case (({drd_req_addr[31:24], drd_req_addr[23:16], drd_req_addr[15:08], drd_req_addr[07:00]} - (base_address_register & 32'hFFFFFFF0)) & 32'hFFFF)
                16'h0000 : rd_rsp_data <= 32'hFEE002F8;
                16'h0010 : rd_rsp_data <= 32'hFEE002F8;
                16'h0020 : rd_rsp_data <= 32'hFEE002F8;
                16'h0030 : rd_rsp_data <= 32'hFEE002F8;
                16'h0040 : rd_rsp_data <= 32'h0020FFFF;
                16'h0044 : rd_rsp_data <= 32'hEBF40004;
                16'h0050 : rd_rsp_data <= 32'h0028FFFF;
                16'h0054 : rd_rsp_data <= 32'hEBF40004;
                16'h0060 : rd_rsp_data <= 32'h0030FFFF;
                16'h0064 : rd_rsp_data <= 32'hEBF40004;
                16'h0070 : rd_rsp_data <= 32'h0038FFFF;
                16'h0074 : rd_rsp_data <= 32'hEBF40004;
                16'h0080 : rd_rsp_data <= 32'h0040FFFF;
                16'h0084 : rd_rsp_data <= 32'hEBF40004;
                16'h0090 : rd_rsp_data <= 32'h0048FFFF;
                16'h0094 : rd_rsp_data <= 32'hEBF40004;
                16'h00A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h00A4 : rd_rsp_data <= 32'hEBF40004;
                16'h00B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h00B4 : rd_rsp_data <= 32'hEBF40004;
                16'h00C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h00C4 : rd_rsp_data <= 32'hEBF40004;
                16'h00D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h00D4 : rd_rsp_data <= 32'hEBF40004;
                16'h00E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h00E4 : rd_rsp_data <= 32'hEBF40004;
                16'h00F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h00F4 : rd_rsp_data <= 32'hEBF40004;
                16'h0104 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0108 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h010C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0110 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0114 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0118 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h011C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0120 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0124 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0128 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h012C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0130 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0134 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0138 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h013C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0140 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0144 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0148 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h014C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0150 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0154 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0158 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h015C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0160 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0164 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0168 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h016C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0170 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0174 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0178 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h017C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0180 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0184 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0188 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h018C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0190 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0194 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0198 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h019C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h01FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0200 : rd_rsp_data <= 32'hFEE002F8;
                16'h0210 : rd_rsp_data <= 32'hFEE002F8;
                16'h0220 : rd_rsp_data <= 32'hFEE002F8;
                16'h0230 : rd_rsp_data <= 32'hFEE002F8;
                16'h0240 : rd_rsp_data <= 32'h0020FFFF;
                16'h0244 : rd_rsp_data <= 32'hEBF40004;
                16'h0250 : rd_rsp_data <= 32'h0028FFFF;
                16'h0254 : rd_rsp_data <= 32'hEBF40004;
                16'h0260 : rd_rsp_data <= 32'h0030FFFF;
                16'h0264 : rd_rsp_data <= 32'hEBF40004;
                16'h0270 : rd_rsp_data <= 32'h0038FFFF;
                16'h0274 : rd_rsp_data <= 32'hEBF40004;
                16'h0280 : rd_rsp_data <= 32'h0040FFFF;
                16'h0284 : rd_rsp_data <= 32'hEBF40004;
                16'h0290 : rd_rsp_data <= 32'h0048FFFF;
                16'h0294 : rd_rsp_data <= 32'hEBF40004;
                16'h02A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h02A4 : rd_rsp_data <= 32'hEBF40004;
                16'h02B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h02B4 : rd_rsp_data <= 32'hEBF40004;
                16'h02C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h02C4 : rd_rsp_data <= 32'hEBF40004;
                16'h02D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h02D4 : rd_rsp_data <= 32'hEBF40004;
                16'h02E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h02E4 : rd_rsp_data <= 32'hEBF40004;
                16'h02F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h02F4 : rd_rsp_data <= 32'hEBF40004;
                16'h0304 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0308 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h030C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0310 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0314 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0318 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h031C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0320 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0324 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0328 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h032C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0330 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0334 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0338 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h033C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0340 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0344 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0348 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h034C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0350 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0354 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0358 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h035C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0360 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0364 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0368 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h036C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0370 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0374 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0378 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h037C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0380 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0384 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0388 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h038C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0390 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0394 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0398 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h039C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h03FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0400 : rd_rsp_data <= 32'hFEE002F8;
                16'h0410 : rd_rsp_data <= 32'hFEE002F8;
                16'h0420 : rd_rsp_data <= 32'hFEE002F8;
                16'h0430 : rd_rsp_data <= 32'hFEE002F8;
                16'h0440 : rd_rsp_data <= 32'h0020FFFF;
                16'h0444 : rd_rsp_data <= 32'hEBF40004;
                16'h0450 : rd_rsp_data <= 32'h0028FFFF;
                16'h0454 : rd_rsp_data <= 32'hEBF40004;
                16'h0460 : rd_rsp_data <= 32'h0030FFFF;
                16'h0464 : rd_rsp_data <= 32'hEBF40004;
                16'h0470 : rd_rsp_data <= 32'h0038FFFF;
                16'h0474 : rd_rsp_data <= 32'hEBF40004;
                16'h0480 : rd_rsp_data <= 32'h0040FFFF;
                16'h0484 : rd_rsp_data <= 32'hEBF40004;
                16'h0490 : rd_rsp_data <= 32'h0048FFFF;
                16'h0494 : rd_rsp_data <= 32'hEBF40004;
                16'h04A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h04A4 : rd_rsp_data <= 32'hEBF40004;
                16'h04B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h04B4 : rd_rsp_data <= 32'hEBF40004;
                16'h04C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h04C4 : rd_rsp_data <= 32'hEBF40004;
                16'h04D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h04D4 : rd_rsp_data <= 32'hEBF40004;
                16'h04E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h04E4 : rd_rsp_data <= 32'hEBF40004;
                16'h04F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h04F4 : rd_rsp_data <= 32'hEBF40004;
                16'h0504 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0508 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h050C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0510 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0514 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0518 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h051C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0520 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0524 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0528 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h052C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0530 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0534 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0538 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h053C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0540 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0544 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0548 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h054C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0550 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0554 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0558 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h055C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0560 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0564 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0568 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h056C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0570 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0574 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0578 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h057C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0580 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0584 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0588 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h058C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0590 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0594 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0598 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h059C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h05FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0600 : rd_rsp_data <= 32'hFEE002F8;
                16'h0610 : rd_rsp_data <= 32'hFEE002F8;
                16'h0620 : rd_rsp_data <= 32'hFEE002F8;
                16'h0630 : rd_rsp_data <= 32'hFEE002F8;
                16'h0640 : rd_rsp_data <= 32'h0020FFFF;
                16'h0644 : rd_rsp_data <= 32'hEBF40004;
                16'h0650 : rd_rsp_data <= 32'h0028FFFF;
                16'h0654 : rd_rsp_data <= 32'hEBF40004;
                16'h0660 : rd_rsp_data <= 32'h0030FFFF;
                16'h0664 : rd_rsp_data <= 32'hEBF40004;
                16'h0670 : rd_rsp_data <= 32'h0038FFFF;
                16'h0674 : rd_rsp_data <= 32'hEBF40004;
                16'h0680 : rd_rsp_data <= 32'h0040FFFF;
                16'h0684 : rd_rsp_data <= 32'hEBF40004;
                16'h0690 : rd_rsp_data <= 32'h0048FFFF;
                16'h0694 : rd_rsp_data <= 32'hEBF40004;
                16'h06A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h06A4 : rd_rsp_data <= 32'hEBF40004;
                16'h06B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h06B4 : rd_rsp_data <= 32'hEBF40004;
                16'h06C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h06C4 : rd_rsp_data <= 32'hEBF40004;
                16'h06D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h06D4 : rd_rsp_data <= 32'hEBF40004;
                16'h06E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h06E4 : rd_rsp_data <= 32'hEBF40004;
                16'h06F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h06F4 : rd_rsp_data <= 32'hEBF40004;
                16'h0704 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0708 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h070C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0710 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0714 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0718 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h071C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0720 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0724 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0728 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h072C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0730 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0734 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0738 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h073C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0740 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0744 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0748 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h074C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0750 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0754 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0758 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h075C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0760 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0764 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0768 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h076C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0770 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0774 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0778 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h077C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0780 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0784 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0788 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h078C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0790 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0794 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0798 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h079C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h07FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0800 : rd_rsp_data <= 32'hFEE002F8;
                16'h0810 : rd_rsp_data <= 32'hFEE002F8;
                16'h0820 : rd_rsp_data <= 32'hFEE002F8;
                16'h0830 : rd_rsp_data <= 32'hFEE002F8;
                16'h0840 : rd_rsp_data <= 32'h0020FFFF;
                16'h0844 : rd_rsp_data <= 32'hEBF40004;
                16'h0850 : rd_rsp_data <= 32'h0028FFFF;
                16'h0854 : rd_rsp_data <= 32'hEBF40004;
                16'h0860 : rd_rsp_data <= 32'h0030FFFF;
                16'h0864 : rd_rsp_data <= 32'hEBF40004;
                16'h0870 : rd_rsp_data <= 32'h0038FFFF;
                16'h0874 : rd_rsp_data <= 32'hEBF40004;
                16'h0880 : rd_rsp_data <= 32'h0040FFFF;
                16'h0884 : rd_rsp_data <= 32'hEBF40004;
                16'h0890 : rd_rsp_data <= 32'h0048FFFF;
                16'h0894 : rd_rsp_data <= 32'hEBF40004;
                16'h08A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h08A4 : rd_rsp_data <= 32'hEBF40004;
                16'h08B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h08B4 : rd_rsp_data <= 32'hEBF40004;
                16'h08C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h08C4 : rd_rsp_data <= 32'hEBF40004;
                16'h08D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h08D4 : rd_rsp_data <= 32'hEBF40004;
                16'h08E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h08E4 : rd_rsp_data <= 32'hEBF40004;
                16'h08F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h08F4 : rd_rsp_data <= 32'hEBF40004;
                16'h0904 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0908 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h090C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0910 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0914 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0918 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h091C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0920 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0924 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0928 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h092C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0930 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0934 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0938 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h093C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0940 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0944 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0948 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h094C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0950 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0954 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0958 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h095C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0960 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0964 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0968 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h096C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0970 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0974 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0978 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h097C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0980 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0984 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0988 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h098C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0990 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0994 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0998 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h099C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h09FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0A00 : rd_rsp_data <= 32'hFEE002F8;
                16'h0A10 : rd_rsp_data <= 32'hFEE002F8;
                16'h0A20 : rd_rsp_data <= 32'hFEE002F8;
                16'h0A30 : rd_rsp_data <= 32'hFEE002F8;
                16'h0A40 : rd_rsp_data <= 32'h0020FFFF;
                16'h0A44 : rd_rsp_data <= 32'hEBF40004;
                16'h0A50 : rd_rsp_data <= 32'h0028FFFF;
                16'h0A54 : rd_rsp_data <= 32'hEBF40004;
                16'h0A60 : rd_rsp_data <= 32'h0030FFFF;
                16'h0A64 : rd_rsp_data <= 32'hEBF40004;
                16'h0A70 : rd_rsp_data <= 32'h0038FFFF;
                16'h0A74 : rd_rsp_data <= 32'hEBF40004;
                16'h0A80 : rd_rsp_data <= 32'h0040FFFF;
                16'h0A84 : rd_rsp_data <= 32'hEBF40004;
                16'h0A90 : rd_rsp_data <= 32'h0048FFFF;
                16'h0A94 : rd_rsp_data <= 32'hEBF40004;
                16'h0AA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h0AA4 : rd_rsp_data <= 32'hEBF40004;
                16'h0AB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h0AB4 : rd_rsp_data <= 32'hEBF40004;
                16'h0AC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h0AC4 : rd_rsp_data <= 32'hEBF40004;
                16'h0AD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h0AD4 : rd_rsp_data <= 32'hEBF40004;
                16'h0AE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h0AE4 : rd_rsp_data <= 32'hEBF40004;
                16'h0AF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h0AF4 : rd_rsp_data <= 32'hEBF40004;
                16'h0B04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0B9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0BFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0C00 : rd_rsp_data <= 32'hFEE002F8;
                16'h0C10 : rd_rsp_data <= 32'hFEE002F8;
                16'h0C20 : rd_rsp_data <= 32'hFEE002F8;
                16'h0C30 : rd_rsp_data <= 32'hFEE002F8;
                16'h0C40 : rd_rsp_data <= 32'h0020FFFF;
                16'h0C44 : rd_rsp_data <= 32'hEBF40004;
                16'h0C50 : rd_rsp_data <= 32'h0028FFFF;
                16'h0C54 : rd_rsp_data <= 32'hEBF40004;
                16'h0C60 : rd_rsp_data <= 32'h0030FFFF;
                16'h0C64 : rd_rsp_data <= 32'hEBF40004;
                16'h0C70 : rd_rsp_data <= 32'h0038FFFF;
                16'h0C74 : rd_rsp_data <= 32'hEBF40004;
                16'h0C80 : rd_rsp_data <= 32'h0040FFFF;
                16'h0C84 : rd_rsp_data <= 32'hEBF40004;
                16'h0C90 : rd_rsp_data <= 32'h0048FFFF;
                16'h0C94 : rd_rsp_data <= 32'hEBF40004;
                16'h0CA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h0CA4 : rd_rsp_data <= 32'hEBF40004;
                16'h0CB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h0CB4 : rd_rsp_data <= 32'hEBF40004;
                16'h0CC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h0CC4 : rd_rsp_data <= 32'hEBF40004;
                16'h0CD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h0CD4 : rd_rsp_data <= 32'hEBF40004;
                16'h0CE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h0CE4 : rd_rsp_data <= 32'hEBF40004;
                16'h0CF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h0CF4 : rd_rsp_data <= 32'hEBF40004;
                16'h0D04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0D9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0DFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0E00 : rd_rsp_data <= 32'hFEE002F8;
                16'h0E10 : rd_rsp_data <= 32'hFEE002F8;
                16'h0E20 : rd_rsp_data <= 32'hFEE002F8;
                16'h0E30 : rd_rsp_data <= 32'hFEE002F8;
                16'h0E40 : rd_rsp_data <= 32'h0020FFFF;
                16'h0E44 : rd_rsp_data <= 32'hEBF40004;
                16'h0E50 : rd_rsp_data <= 32'h0028FFFF;
                16'h0E54 : rd_rsp_data <= 32'hEBF40004;
                16'h0E60 : rd_rsp_data <= 32'h0030FFFF;
                16'h0E64 : rd_rsp_data <= 32'hEBF40004;
                16'h0E70 : rd_rsp_data <= 32'h0038FFFF;
                16'h0E74 : rd_rsp_data <= 32'hEBF40004;
                16'h0E80 : rd_rsp_data <= 32'h0040FFFF;
                16'h0E84 : rd_rsp_data <= 32'hEBF40004;
                16'h0E90 : rd_rsp_data <= 32'h0048FFFF;
                16'h0E94 : rd_rsp_data <= 32'hEBF40004;
                16'h0EA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h0EA4 : rd_rsp_data <= 32'hEBF40004;
                16'h0EB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h0EB4 : rd_rsp_data <= 32'hEBF40004;
                16'h0EC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h0EC4 : rd_rsp_data <= 32'hEBF40004;
                16'h0ED0 : rd_rsp_data <= 32'h0068FFFF;
                16'h0ED4 : rd_rsp_data <= 32'hEBF40004;
                16'h0EE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h0EE4 : rd_rsp_data <= 32'hEBF40004;
                16'h0EF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h0EF4 : rd_rsp_data <= 32'hEBF40004;
                16'h0F04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0F9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0FFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1000 : rd_rsp_data <= 32'hFEE002F8;
                16'h1010 : rd_rsp_data <= 32'hFEE002F8;
                16'h1020 : rd_rsp_data <= 32'hFEE002F8;
                16'h1030 : rd_rsp_data <= 32'hFEE002F8;
                16'h1040 : rd_rsp_data <= 32'h0020FFFF;
                16'h1044 : rd_rsp_data <= 32'hEBF40004;
                16'h1050 : rd_rsp_data <= 32'h0028FFFF;
                16'h1054 : rd_rsp_data <= 32'hEBF40004;
                16'h1060 : rd_rsp_data <= 32'h0030FFFF;
                16'h1064 : rd_rsp_data <= 32'hEBF40004;
                16'h1070 : rd_rsp_data <= 32'h0038FFFF;
                16'h1074 : rd_rsp_data <= 32'hEBF40004;
                16'h1080 : rd_rsp_data <= 32'h0040FFFF;
                16'h1084 : rd_rsp_data <= 32'hEBF40004;
                16'h1090 : rd_rsp_data <= 32'h0048FFFF;
                16'h1094 : rd_rsp_data <= 32'hEBF40004;
                16'h10A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h10A4 : rd_rsp_data <= 32'hEBF40004;
                16'h10B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h10B4 : rd_rsp_data <= 32'hEBF40004;
                16'h10C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h10C4 : rd_rsp_data <= 32'hEBF40004;
                16'h10D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h10D4 : rd_rsp_data <= 32'hEBF40004;
                16'h10E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h10E4 : rd_rsp_data <= 32'hEBF40004;
                16'h10F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h10F4 : rd_rsp_data <= 32'hEBF40004;
                16'h1104 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1108 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h110C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1110 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1114 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1118 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h111C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1120 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1124 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1128 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h112C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1130 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1134 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1138 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h113C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1140 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1144 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1148 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h114C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1150 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1154 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1158 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h115C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1160 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1164 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1168 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h116C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1170 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1174 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1178 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h117C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1180 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1184 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1188 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h118C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1190 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1194 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1198 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h119C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h11FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1200 : rd_rsp_data <= 32'hFEE002F8;
                16'h1210 : rd_rsp_data <= 32'hFEE002F8;
                16'h1220 : rd_rsp_data <= 32'hFEE002F8;
                16'h1230 : rd_rsp_data <= 32'hFEE002F8;
                16'h1240 : rd_rsp_data <= 32'h0020FFFF;
                16'h1244 : rd_rsp_data <= 32'hEBF40004;
                16'h1250 : rd_rsp_data <= 32'h0028FFFF;
                16'h1254 : rd_rsp_data <= 32'hEBF40004;
                16'h1260 : rd_rsp_data <= 32'h0030FFFF;
                16'h1264 : rd_rsp_data <= 32'hEBF40004;
                16'h1270 : rd_rsp_data <= 32'h0038FFFF;
                16'h1274 : rd_rsp_data <= 32'hEBF40004;
                16'h1280 : rd_rsp_data <= 32'h0040FFFF;
                16'h1284 : rd_rsp_data <= 32'hEBF40004;
                16'h1290 : rd_rsp_data <= 32'h0048FFFF;
                16'h1294 : rd_rsp_data <= 32'hEBF40004;
                16'h12A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h12A4 : rd_rsp_data <= 32'hEBF40004;
                16'h12B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h12B4 : rd_rsp_data <= 32'hEBF40004;
                16'h12C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h12C4 : rd_rsp_data <= 32'hEBF40004;
                16'h12D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h12D4 : rd_rsp_data <= 32'hEBF40004;
                16'h12E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h12E4 : rd_rsp_data <= 32'hEBF40004;
                16'h12F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h12F4 : rd_rsp_data <= 32'hEBF40004;
                16'h1304 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1308 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h130C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1310 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1314 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1318 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h131C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1320 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1324 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1328 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h132C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1330 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1334 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1338 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h133C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1340 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1344 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1348 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h134C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1350 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1354 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1358 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h135C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1360 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1364 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1368 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h136C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1370 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1374 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1378 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h137C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1380 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1384 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1388 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h138C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1390 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1394 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1398 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h139C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h13FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1400 : rd_rsp_data <= 32'hFEE002F8;
                16'h1410 : rd_rsp_data <= 32'hFEE002F8;
                16'h1420 : rd_rsp_data <= 32'hFEE002F8;
                16'h1430 : rd_rsp_data <= 32'hFEE002F8;
                16'h1440 : rd_rsp_data <= 32'h0020FFFF;
                16'h1444 : rd_rsp_data <= 32'hEBF40004;
                16'h1450 : rd_rsp_data <= 32'h0028FFFF;
                16'h1454 : rd_rsp_data <= 32'hEBF40004;
                16'h1460 : rd_rsp_data <= 32'h0030FFFF;
                16'h1464 : rd_rsp_data <= 32'hEBF40004;
                16'h1470 : rd_rsp_data <= 32'h0038FFFF;
                16'h1474 : rd_rsp_data <= 32'hEBF40004;
                16'h1480 : rd_rsp_data <= 32'h0040FFFF;
                16'h1484 : rd_rsp_data <= 32'hEBF40004;
                16'h1490 : rd_rsp_data <= 32'h0048FFFF;
                16'h1494 : rd_rsp_data <= 32'hEBF40004;
                16'h14A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h14A4 : rd_rsp_data <= 32'hEBF40004;
                16'h14B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h14B4 : rd_rsp_data <= 32'hEBF40004;
                16'h14C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h14C4 : rd_rsp_data <= 32'hEBF40004;
                16'h14D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h14D4 : rd_rsp_data <= 32'hEBF40004;
                16'h14E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h14E4 : rd_rsp_data <= 32'hEBF40004;
                16'h14F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h14F4 : rd_rsp_data <= 32'hEBF40004;
                16'h1504 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1508 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h150C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1510 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1514 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1518 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h151C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1520 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1524 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1528 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h152C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1530 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1534 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1538 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h153C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1540 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1544 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1548 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h154C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1550 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1554 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1558 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h155C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1560 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1564 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1568 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h156C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1570 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1574 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1578 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h157C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1580 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1584 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1588 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h158C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1590 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1594 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1598 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h159C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h15FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1600 : rd_rsp_data <= 32'hFEE002F8;
                16'h1610 : rd_rsp_data <= 32'hFEE002F8;
                16'h1620 : rd_rsp_data <= 32'hFEE002F8;
                16'h1630 : rd_rsp_data <= 32'hFEE002F8;
                16'h1640 : rd_rsp_data <= 32'h0020FFFF;
                16'h1644 : rd_rsp_data <= 32'hEBF40004;
                16'h1650 : rd_rsp_data <= 32'h0028FFFF;
                16'h1654 : rd_rsp_data <= 32'hEBF40004;
                16'h1660 : rd_rsp_data <= 32'h0030FFFF;
                16'h1664 : rd_rsp_data <= 32'hEBF40004;
                16'h1670 : rd_rsp_data <= 32'h0038FFFF;
                16'h1674 : rd_rsp_data <= 32'hEBF40004;
                16'h1680 : rd_rsp_data <= 32'h0040FFFF;
                16'h1684 : rd_rsp_data <= 32'hEBF40004;
                16'h1690 : rd_rsp_data <= 32'h0048FFFF;
                16'h1694 : rd_rsp_data <= 32'hEBF40004;
                16'h16A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h16A4 : rd_rsp_data <= 32'hEBF40004;
                16'h16B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h16B4 : rd_rsp_data <= 32'hEBF40004;
                16'h16C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h16C4 : rd_rsp_data <= 32'hEBF40004;
                16'h16D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h16D4 : rd_rsp_data <= 32'hEBF40004;
                16'h16E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h16E4 : rd_rsp_data <= 32'hEBF40004;
                16'h16F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h16F4 : rd_rsp_data <= 32'hEBF40004;
                16'h1704 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1708 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h170C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1710 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1714 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1718 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h171C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1720 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1724 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1728 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h172C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1730 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1734 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1738 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h173C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1740 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1744 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1748 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h174C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1750 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1754 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1758 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h175C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1760 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1764 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1768 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h176C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1770 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1774 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1778 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h177C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1780 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1784 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1788 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h178C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1790 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1794 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1798 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h179C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h17FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1800 : rd_rsp_data <= 32'hFEE002F8;
                16'h1810 : rd_rsp_data <= 32'hFEE002F8;
                16'h1820 : rd_rsp_data <= 32'hFEE002F8;
                16'h1830 : rd_rsp_data <= 32'hFEE002F8;
                16'h1840 : rd_rsp_data <= 32'h0020FFFF;
                16'h1844 : rd_rsp_data <= 32'hEBF40004;
                16'h1850 : rd_rsp_data <= 32'h0028FFFF;
                16'h1854 : rd_rsp_data <= 32'hEBF40004;
                16'h1860 : rd_rsp_data <= 32'h0030FFFF;
                16'h1864 : rd_rsp_data <= 32'hEBF40004;
                16'h1870 : rd_rsp_data <= 32'h0038FFFF;
                16'h1874 : rd_rsp_data <= 32'hEBF40004;
                16'h1880 : rd_rsp_data <= 32'h0040FFFF;
                16'h1884 : rd_rsp_data <= 32'hEBF40004;
                16'h1890 : rd_rsp_data <= 32'h0048FFFF;
                16'h1894 : rd_rsp_data <= 32'hEBF40004;
                16'h18A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h18A4 : rd_rsp_data <= 32'hEBF40004;
                16'h18B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h18B4 : rd_rsp_data <= 32'hEBF40004;
                16'h18C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h18C4 : rd_rsp_data <= 32'hEBF40004;
                16'h18D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h18D4 : rd_rsp_data <= 32'hEBF40004;
                16'h18E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h18E4 : rd_rsp_data <= 32'hEBF40004;
                16'h18F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h18F4 : rd_rsp_data <= 32'hEBF40004;
                16'h1904 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1908 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h190C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1910 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1914 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1918 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h191C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1920 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1924 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1928 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h192C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1930 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1934 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1938 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h193C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1940 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1944 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1948 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h194C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1950 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1954 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1958 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h195C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1960 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1964 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1968 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h196C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1970 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1974 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1978 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h197C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1980 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1984 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1988 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h198C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1990 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1994 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1998 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h199C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h19FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1A00 : rd_rsp_data <= 32'hFEE002F8;
                16'h1A10 : rd_rsp_data <= 32'hFEE002F8;
                16'h1A20 : rd_rsp_data <= 32'hFEE002F8;
                16'h1A30 : rd_rsp_data <= 32'hFEE002F8;
                16'h1A40 : rd_rsp_data <= 32'h0020FFFF;
                16'h1A44 : rd_rsp_data <= 32'hEBF40004;
                16'h1A50 : rd_rsp_data <= 32'h0028FFFF;
                16'h1A54 : rd_rsp_data <= 32'hEBF40004;
                16'h1A60 : rd_rsp_data <= 32'h0030FFFF;
                16'h1A64 : rd_rsp_data <= 32'hEBF40004;
                16'h1A70 : rd_rsp_data <= 32'h0038FFFF;
                16'h1A74 : rd_rsp_data <= 32'hEBF40004;
                16'h1A80 : rd_rsp_data <= 32'h0040FFFF;
                16'h1A84 : rd_rsp_data <= 32'hEBF40004;
                16'h1A90 : rd_rsp_data <= 32'h0048FFFF;
                16'h1A94 : rd_rsp_data <= 32'hEBF40004;
                16'h1AA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h1AA4 : rd_rsp_data <= 32'hEBF40004;
                16'h1AB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h1AB4 : rd_rsp_data <= 32'hEBF40004;
                16'h1AC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h1AC4 : rd_rsp_data <= 32'hEBF40004;
                16'h1AD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h1AD4 : rd_rsp_data <= 32'hEBF40004;
                16'h1AE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h1AE4 : rd_rsp_data <= 32'hEBF40004;
                16'h1AF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h1AF4 : rd_rsp_data <= 32'hEBF40004;
                16'h1B04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1B9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1BFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1C00 : rd_rsp_data <= 32'hFEE002F8;
                16'h1C10 : rd_rsp_data <= 32'hFEE002F8;
                16'h1C20 : rd_rsp_data <= 32'hFEE002F8;
                16'h1C30 : rd_rsp_data <= 32'hFEE002F8;
                16'h1C40 : rd_rsp_data <= 32'h0020FFFF;
                16'h1C44 : rd_rsp_data <= 32'hEBF40004;
                16'h1C50 : rd_rsp_data <= 32'h0028FFFF;
                16'h1C54 : rd_rsp_data <= 32'hEBF40004;
                16'h1C60 : rd_rsp_data <= 32'h0030FFFF;
                16'h1C64 : rd_rsp_data <= 32'hEBF40004;
                16'h1C70 : rd_rsp_data <= 32'h0038FFFF;
                16'h1C74 : rd_rsp_data <= 32'hEBF40004;
                16'h1C80 : rd_rsp_data <= 32'h0040FFFF;
                16'h1C84 : rd_rsp_data <= 32'hEBF40004;
                16'h1C90 : rd_rsp_data <= 32'h0048FFFF;
                16'h1C94 : rd_rsp_data <= 32'hEBF40004;
                16'h1CA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h1CA4 : rd_rsp_data <= 32'hEBF40004;
                16'h1CB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h1CB4 : rd_rsp_data <= 32'hEBF40004;
                16'h1CC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h1CC4 : rd_rsp_data <= 32'hEBF40004;
                16'h1CD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h1CD4 : rd_rsp_data <= 32'hEBF40004;
                16'h1CE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h1CE4 : rd_rsp_data <= 32'hEBF40004;
                16'h1CF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h1CF4 : rd_rsp_data <= 32'hEBF40004;
                16'h1D04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1D9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1DFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1E00 : rd_rsp_data <= 32'hFEE002F8;
                16'h1E10 : rd_rsp_data <= 32'hFEE002F8;
                16'h1E20 : rd_rsp_data <= 32'hFEE002F8;
                16'h1E30 : rd_rsp_data <= 32'hFEE002F8;
                16'h1E40 : rd_rsp_data <= 32'h0020FFFF;
                16'h1E44 : rd_rsp_data <= 32'hEBF40004;
                16'h1E50 : rd_rsp_data <= 32'h0028FFFF;
                16'h1E54 : rd_rsp_data <= 32'hEBF40004;
                16'h1E60 : rd_rsp_data <= 32'h0030FFFF;
                16'h1E64 : rd_rsp_data <= 32'hEBF40004;
                16'h1E70 : rd_rsp_data <= 32'h0038FFFF;
                16'h1E74 : rd_rsp_data <= 32'hEBF40004;
                16'h1E80 : rd_rsp_data <= 32'h0040FFFF;
                16'h1E84 : rd_rsp_data <= 32'hEBF40004;
                16'h1E90 : rd_rsp_data <= 32'h0048FFFF;
                16'h1E94 : rd_rsp_data <= 32'hEBF40004;
                16'h1EA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h1EA4 : rd_rsp_data <= 32'hEBF40004;
                16'h1EB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h1EB4 : rd_rsp_data <= 32'hEBF40004;
                16'h1EC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h1EC4 : rd_rsp_data <= 32'hEBF40004;
                16'h1ED0 : rd_rsp_data <= 32'h0068FFFF;
                16'h1ED4 : rd_rsp_data <= 32'hEBF40004;
                16'h1EE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h1EE4 : rd_rsp_data <= 32'hEBF40004;
                16'h1EF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h1EF4 : rd_rsp_data <= 32'hEBF40004;
                16'h1F04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1F9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h1FFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2000 : rd_rsp_data <= 32'hFEE002F8;
                16'h2010 : rd_rsp_data <= 32'hFEE002F8;
                16'h2020 : rd_rsp_data <= 32'hFEE002F8;
                16'h2030 : rd_rsp_data <= 32'hFEE002F8;
                16'h2040 : rd_rsp_data <= 32'h0020FFFF;
                16'h2044 : rd_rsp_data <= 32'hEBF40004;
                16'h2050 : rd_rsp_data <= 32'h0028FFFF;
                16'h2054 : rd_rsp_data <= 32'hEBF40004;
                16'h2060 : rd_rsp_data <= 32'h0030FFFF;
                16'h2064 : rd_rsp_data <= 32'hEBF40004;
                16'h2070 : rd_rsp_data <= 32'h0038FFFF;
                16'h2074 : rd_rsp_data <= 32'hEBF40004;
                16'h2080 : rd_rsp_data <= 32'h0040FFFF;
                16'h2084 : rd_rsp_data <= 32'hEBF40004;
                16'h2090 : rd_rsp_data <= 32'h0048FFFF;
                16'h2094 : rd_rsp_data <= 32'hEBF40004;
                16'h20A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h20A4 : rd_rsp_data <= 32'hEBF40004;
                16'h20B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h20B4 : rd_rsp_data <= 32'hEBF40004;
                16'h20C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h20C4 : rd_rsp_data <= 32'hEBF40004;
                16'h20D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h20D4 : rd_rsp_data <= 32'hEBF40004;
                16'h20E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h20E4 : rd_rsp_data <= 32'hEBF40004;
                16'h20F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h20F4 : rd_rsp_data <= 32'hEBF40004;
                16'h2104 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2108 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h210C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2110 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2114 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2118 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h211C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2120 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2124 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2128 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h212C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2130 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2134 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2138 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h213C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2140 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2144 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2148 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h214C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2150 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2154 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2158 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h215C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2160 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2164 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2168 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h216C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2170 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2174 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2178 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h217C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2180 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2184 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2188 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h218C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2190 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2194 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2198 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h219C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h21FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2200 : rd_rsp_data <= 32'hFEE002F8;
                16'h2210 : rd_rsp_data <= 32'hFEE002F8;
                16'h2220 : rd_rsp_data <= 32'hFEE002F8;
                16'h2230 : rd_rsp_data <= 32'hFEE002F8;
                16'h2240 : rd_rsp_data <= 32'h0020FFFF;
                16'h2244 : rd_rsp_data <= 32'hEBF40004;
                16'h2250 : rd_rsp_data <= 32'h0028FFFF;
                16'h2254 : rd_rsp_data <= 32'hEBF40004;
                16'h2260 : rd_rsp_data <= 32'h0030FFFF;
                16'h2264 : rd_rsp_data <= 32'hEBF40004;
                16'h2270 : rd_rsp_data <= 32'h0038FFFF;
                16'h2274 : rd_rsp_data <= 32'hEBF40004;
                16'h2280 : rd_rsp_data <= 32'h0040FFFF;
                16'h2284 : rd_rsp_data <= 32'hEBF40004;
                16'h2290 : rd_rsp_data <= 32'h0048FFFF;
                16'h2294 : rd_rsp_data <= 32'hEBF40004;
                16'h22A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h22A4 : rd_rsp_data <= 32'hEBF40004;
                16'h22B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h22B4 : rd_rsp_data <= 32'hEBF40004;
                16'h22C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h22C4 : rd_rsp_data <= 32'hEBF40004;
                16'h22D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h22D4 : rd_rsp_data <= 32'hEBF40004;
                16'h22E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h22E4 : rd_rsp_data <= 32'hEBF40004;
                16'h22F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h22F4 : rd_rsp_data <= 32'hEBF40004;
                16'h2304 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2308 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h230C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2310 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2314 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2318 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h231C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2320 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2324 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2328 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h232C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2330 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2334 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2338 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h233C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2340 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2344 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2348 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h234C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2350 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2354 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2358 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h235C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2360 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2364 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2368 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h236C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2370 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2374 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2378 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h237C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2380 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2384 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2388 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h238C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2390 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2394 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2398 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h239C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h23FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2400 : rd_rsp_data <= 32'hFEE002F8;
                16'h2410 : rd_rsp_data <= 32'hFEE002F8;
                16'h2420 : rd_rsp_data <= 32'hFEE002F8;
                16'h2430 : rd_rsp_data <= 32'hFEE002F8;
                16'h2440 : rd_rsp_data <= 32'h0020FFFF;
                16'h2444 : rd_rsp_data <= 32'hEBF40004;
                16'h2450 : rd_rsp_data <= 32'h0028FFFF;
                16'h2454 : rd_rsp_data <= 32'hEBF40004;
                16'h2460 : rd_rsp_data <= 32'h0030FFFF;
                16'h2464 : rd_rsp_data <= 32'hEBF40004;
                16'h2470 : rd_rsp_data <= 32'h0038FFFF;
                16'h2474 : rd_rsp_data <= 32'hEBF40004;
                16'h2480 : rd_rsp_data <= 32'h0040FFFF;
                16'h2484 : rd_rsp_data <= 32'hEBF40004;
                16'h2490 : rd_rsp_data <= 32'h0048FFFF;
                16'h2494 : rd_rsp_data <= 32'hEBF40004;
                16'h24A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h24A4 : rd_rsp_data <= 32'hEBF40004;
                16'h24B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h24B4 : rd_rsp_data <= 32'hEBF40004;
                16'h24C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h24C4 : rd_rsp_data <= 32'hEBF40004;
                16'h24D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h24D4 : rd_rsp_data <= 32'hEBF40004;
                16'h24E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h24E4 : rd_rsp_data <= 32'hEBF40004;
                16'h24F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h24F4 : rd_rsp_data <= 32'hEBF40004;
                16'h2504 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2508 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h250C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2510 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2514 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2518 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h251C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2520 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2524 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2528 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h252C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2530 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2534 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2538 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h253C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2540 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2544 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2548 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h254C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2550 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2554 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2558 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h255C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2560 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2564 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2568 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h256C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2570 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2574 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2578 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h257C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2580 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2584 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2588 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h258C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2590 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2594 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2598 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h259C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h25FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2600 : rd_rsp_data <= 32'hFEE002F8;
                16'h2610 : rd_rsp_data <= 32'hFEE002F8;
                16'h2620 : rd_rsp_data <= 32'hFEE002F8;
                16'h2630 : rd_rsp_data <= 32'hFEE002F8;
                16'h2640 : rd_rsp_data <= 32'h0020FFFF;
                16'h2644 : rd_rsp_data <= 32'hEBF40004;
                16'h2650 : rd_rsp_data <= 32'h0028FFFF;
                16'h2654 : rd_rsp_data <= 32'hEBF40004;
                16'h2660 : rd_rsp_data <= 32'h0030FFFF;
                16'h2664 : rd_rsp_data <= 32'hEBF40004;
                16'h2670 : rd_rsp_data <= 32'h0038FFFF;
                16'h2674 : rd_rsp_data <= 32'hEBF40004;
                16'h2680 : rd_rsp_data <= 32'h0040FFFF;
                16'h2684 : rd_rsp_data <= 32'hEBF40004;
                16'h2690 : rd_rsp_data <= 32'h0048FFFF;
                16'h2694 : rd_rsp_data <= 32'hEBF40004;
                16'h26A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h26A4 : rd_rsp_data <= 32'hEBF40004;
                16'h26B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h26B4 : rd_rsp_data <= 32'hEBF40004;
                16'h26C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h26C4 : rd_rsp_data <= 32'hEBF40004;
                16'h26D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h26D4 : rd_rsp_data <= 32'hEBF40004;
                16'h26E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h26E4 : rd_rsp_data <= 32'hEBF40004;
                16'h26F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h26F4 : rd_rsp_data <= 32'hEBF40004;
                16'h2704 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2708 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h270C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2710 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2714 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2718 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h271C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2720 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2724 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2728 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h272C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2730 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2734 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2738 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h273C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2740 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2744 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2748 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h274C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2750 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2754 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2758 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h275C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2760 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2764 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2768 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h276C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2770 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2774 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2778 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h277C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2780 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2784 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2788 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h278C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2790 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2794 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2798 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h279C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h27FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2800 : rd_rsp_data <= 32'hFEE002F8;
                16'h2810 : rd_rsp_data <= 32'hFEE002F8;
                16'h2820 : rd_rsp_data <= 32'hFEE002F8;
                16'h2830 : rd_rsp_data <= 32'hFEE002F8;
                16'h2840 : rd_rsp_data <= 32'h0020FFFF;
                16'h2844 : rd_rsp_data <= 32'hEBF40004;
                16'h2850 : rd_rsp_data <= 32'h0028FFFF;
                16'h2854 : rd_rsp_data <= 32'hEBF40004;
                16'h2860 : rd_rsp_data <= 32'h0030FFFF;
                16'h2864 : rd_rsp_data <= 32'hEBF40004;
                16'h2870 : rd_rsp_data <= 32'h0038FFFF;
                16'h2874 : rd_rsp_data <= 32'hEBF40004;
                16'h2880 : rd_rsp_data <= 32'h0040FFFF;
                16'h2884 : rd_rsp_data <= 32'hEBF40004;
                16'h2890 : rd_rsp_data <= 32'h0048FFFF;
                16'h2894 : rd_rsp_data <= 32'hEBF40004;
                16'h28A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h28A4 : rd_rsp_data <= 32'hEBF40004;
                16'h28B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h28B4 : rd_rsp_data <= 32'hEBF40004;
                16'h28C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h28C4 : rd_rsp_data <= 32'hEBF40004;
                16'h28D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h28D4 : rd_rsp_data <= 32'hEBF40004;
                16'h28E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h28E4 : rd_rsp_data <= 32'hEBF40004;
                16'h28F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h28F4 : rd_rsp_data <= 32'hEBF40004;
                16'h2904 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2908 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h290C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2910 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2914 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2918 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h291C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2920 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2924 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2928 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h292C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2930 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2934 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2938 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h293C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2940 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2944 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2948 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h294C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2950 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2954 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2958 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h295C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2960 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2964 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2968 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h296C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2970 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2974 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2978 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h297C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2980 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2984 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2988 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h298C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2990 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2994 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2998 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h299C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h29FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2A00 : rd_rsp_data <= 32'hFEE002F8;
                16'h2A10 : rd_rsp_data <= 32'hFEE002F8;
                16'h2A20 : rd_rsp_data <= 32'hFEE002F8;
                16'h2A30 : rd_rsp_data <= 32'hFEE002F8;
                16'h2A40 : rd_rsp_data <= 32'h0020FFFF;
                16'h2A44 : rd_rsp_data <= 32'hEBF40004;
                16'h2A50 : rd_rsp_data <= 32'h0028FFFF;
                16'h2A54 : rd_rsp_data <= 32'hEBF40004;
                16'h2A60 : rd_rsp_data <= 32'h0030FFFF;
                16'h2A64 : rd_rsp_data <= 32'hEBF40004;
                16'h2A70 : rd_rsp_data <= 32'h0038FFFF;
                16'h2A74 : rd_rsp_data <= 32'hEBF40004;
                16'h2A80 : rd_rsp_data <= 32'h0040FFFF;
                16'h2A84 : rd_rsp_data <= 32'hEBF40004;
                16'h2A90 : rd_rsp_data <= 32'h0048FFFF;
                16'h2A94 : rd_rsp_data <= 32'hEBF40004;
                16'h2AA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h2AA4 : rd_rsp_data <= 32'hEBF40004;
                16'h2AB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h2AB4 : rd_rsp_data <= 32'hEBF40004;
                16'h2AC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h2AC4 : rd_rsp_data <= 32'hEBF40004;
                16'h2AD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h2AD4 : rd_rsp_data <= 32'hEBF40004;
                16'h2AE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h2AE4 : rd_rsp_data <= 32'hEBF40004;
                16'h2AF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h2AF4 : rd_rsp_data <= 32'hEBF40004;
                16'h2B04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2B9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2BFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2C00 : rd_rsp_data <= 32'hFEE002F8;
                16'h2C10 : rd_rsp_data <= 32'hFEE002F8;
                16'h2C20 : rd_rsp_data <= 32'hFEE002F8;
                16'h2C30 : rd_rsp_data <= 32'hFEE002F8;
                16'h2C40 : rd_rsp_data <= 32'h0020FFFF;
                16'h2C44 : rd_rsp_data <= 32'hEBF40004;
                16'h2C50 : rd_rsp_data <= 32'h0028FFFF;
                16'h2C54 : rd_rsp_data <= 32'hEBF40004;
                16'h2C60 : rd_rsp_data <= 32'h0030FFFF;
                16'h2C64 : rd_rsp_data <= 32'hEBF40004;
                16'h2C70 : rd_rsp_data <= 32'h0038FFFF;
                16'h2C74 : rd_rsp_data <= 32'hEBF40004;
                16'h2C80 : rd_rsp_data <= 32'h0040FFFF;
                16'h2C84 : rd_rsp_data <= 32'hEBF40004;
                16'h2C90 : rd_rsp_data <= 32'h0048FFFF;
                16'h2C94 : rd_rsp_data <= 32'hEBF40004;
                16'h2CA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h2CA4 : rd_rsp_data <= 32'hEBF40004;
                16'h2CB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h2CB4 : rd_rsp_data <= 32'hEBF40004;
                16'h2CC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h2CC4 : rd_rsp_data <= 32'hEBF40004;
                16'h2CD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h2CD4 : rd_rsp_data <= 32'hEBF40004;
                16'h2CE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h2CE4 : rd_rsp_data <= 32'hEBF40004;
                16'h2CF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h2CF4 : rd_rsp_data <= 32'hEBF40004;
                16'h2D04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2D9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2DFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2E00 : rd_rsp_data <= 32'hFEE002F8;
                16'h2E10 : rd_rsp_data <= 32'hFEE002F8;
                16'h2E20 : rd_rsp_data <= 32'hFEE002F8;
                16'h2E30 : rd_rsp_data <= 32'hFEE002F8;
                16'h2E40 : rd_rsp_data <= 32'h0020FFFF;
                16'h2E44 : rd_rsp_data <= 32'hEBF40004;
                16'h2E50 : rd_rsp_data <= 32'h0028FFFF;
                16'h2E54 : rd_rsp_data <= 32'hEBF40004;
                16'h2E60 : rd_rsp_data <= 32'h0030FFFF;
                16'h2E64 : rd_rsp_data <= 32'hEBF40004;
                16'h2E70 : rd_rsp_data <= 32'h0038FFFF;
                16'h2E74 : rd_rsp_data <= 32'hEBF40004;
                16'h2E80 : rd_rsp_data <= 32'h0040FFFF;
                16'h2E84 : rd_rsp_data <= 32'hEBF40004;
                16'h2E90 : rd_rsp_data <= 32'h0048FFFF;
                16'h2E94 : rd_rsp_data <= 32'hEBF40004;
                16'h2EA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h2EA4 : rd_rsp_data <= 32'hEBF40004;
                16'h2EB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h2EB4 : rd_rsp_data <= 32'hEBF40004;
                16'h2EC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h2EC4 : rd_rsp_data <= 32'hEBF40004;
                16'h2ED0 : rd_rsp_data <= 32'h0068FFFF;
                16'h2ED4 : rd_rsp_data <= 32'hEBF40004;
                16'h2EE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h2EE4 : rd_rsp_data <= 32'hEBF40004;
                16'h2EF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h2EF4 : rd_rsp_data <= 32'hEBF40004;
                16'h2F04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2F9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h2FFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3000 : rd_rsp_data <= 32'hFEE002F8;
                16'h3010 : rd_rsp_data <= 32'hFEE002F8;
                16'h3020 : rd_rsp_data <= 32'hFEE002F8;
                16'h3030 : rd_rsp_data <= 32'hFEE002F8;
                16'h3040 : rd_rsp_data <= 32'h0020FFFF;
                16'h3044 : rd_rsp_data <= 32'hEBF40004;
                16'h3050 : rd_rsp_data <= 32'h0028FFFF;
                16'h3054 : rd_rsp_data <= 32'hEBF40004;
                16'h3060 : rd_rsp_data <= 32'h0030FFFF;
                16'h3064 : rd_rsp_data <= 32'hEBF40004;
                16'h3070 : rd_rsp_data <= 32'h0038FFFF;
                16'h3074 : rd_rsp_data <= 32'hEBF40004;
                16'h3080 : rd_rsp_data <= 32'h0040FFFF;
                16'h3084 : rd_rsp_data <= 32'hEBF40004;
                16'h3090 : rd_rsp_data <= 32'h0048FFFF;
                16'h3094 : rd_rsp_data <= 32'hEBF40004;
                16'h30A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h30A4 : rd_rsp_data <= 32'hEBF40004;
                16'h30B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h30B4 : rd_rsp_data <= 32'hEBF40004;
                16'h30C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h30C4 : rd_rsp_data <= 32'hEBF40004;
                16'h30D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h30D4 : rd_rsp_data <= 32'hEBF40004;
                16'h30E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h30E4 : rd_rsp_data <= 32'hEBF40004;
                16'h30F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h30F4 : rd_rsp_data <= 32'hEBF40004;
                16'h3104 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3108 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h310C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3110 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3114 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3118 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h311C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3120 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3124 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3128 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h312C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3130 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3134 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3138 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h313C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3140 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3144 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3148 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h314C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3150 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3154 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3158 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h315C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3160 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3164 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3168 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h316C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3170 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3174 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3178 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h317C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3180 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3184 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3188 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h318C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3190 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3194 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3198 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h319C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h31FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3200 : rd_rsp_data <= 32'hFEE002F8;
                16'h3210 : rd_rsp_data <= 32'hFEE002F8;
                16'h3220 : rd_rsp_data <= 32'hFEE002F8;
                16'h3230 : rd_rsp_data <= 32'hFEE002F8;
                16'h3240 : rd_rsp_data <= 32'h0020FFFF;
                16'h3244 : rd_rsp_data <= 32'hEBF40004;
                16'h3250 : rd_rsp_data <= 32'h0028FFFF;
                16'h3254 : rd_rsp_data <= 32'hEBF40004;
                16'h3260 : rd_rsp_data <= 32'h0030FFFF;
                16'h3264 : rd_rsp_data <= 32'hEBF40004;
                16'h3270 : rd_rsp_data <= 32'h0038FFFF;
                16'h3274 : rd_rsp_data <= 32'hEBF40004;
                16'h3280 : rd_rsp_data <= 32'h0040FFFF;
                16'h3284 : rd_rsp_data <= 32'hEBF40004;
                16'h3290 : rd_rsp_data <= 32'h0048FFFF;
                16'h3294 : rd_rsp_data <= 32'hEBF40004;
                16'h32A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h32A4 : rd_rsp_data <= 32'hEBF40004;
                16'h32B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h32B4 : rd_rsp_data <= 32'hEBF40004;
                16'h32C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h32C4 : rd_rsp_data <= 32'hEBF40004;
                16'h32D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h32D4 : rd_rsp_data <= 32'hEBF40004;
                16'h32E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h32E4 : rd_rsp_data <= 32'hEBF40004;
                16'h32F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h32F4 : rd_rsp_data <= 32'hEBF40004;
                16'h3304 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3308 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h330C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3310 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3314 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3318 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h331C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3320 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3324 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3328 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h332C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3330 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3334 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3338 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h333C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3340 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3344 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3348 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h334C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3350 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3354 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3358 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h335C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3360 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3364 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3368 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h336C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3370 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3374 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3378 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h337C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3380 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3384 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3388 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h338C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3390 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3394 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3398 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h339C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h33FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3400 : rd_rsp_data <= 32'hFEE002F8;
                16'h3410 : rd_rsp_data <= 32'hFEE002F8;
                16'h3420 : rd_rsp_data <= 32'hFEE002F8;
                16'h3430 : rd_rsp_data <= 32'hFEE002F8;
                16'h3440 : rd_rsp_data <= 32'h0020FFFF;
                16'h3444 : rd_rsp_data <= 32'hEBF40004;
                16'h3450 : rd_rsp_data <= 32'h0028FFFF;
                16'h3454 : rd_rsp_data <= 32'hEBF40004;
                16'h3460 : rd_rsp_data <= 32'h0030FFFF;
                16'h3464 : rd_rsp_data <= 32'hEBF40004;
                16'h3470 : rd_rsp_data <= 32'h0038FFFF;
                16'h3474 : rd_rsp_data <= 32'hEBF40004;
                16'h3480 : rd_rsp_data <= 32'h0040FFFF;
                16'h3484 : rd_rsp_data <= 32'hEBF40004;
                16'h3490 : rd_rsp_data <= 32'h0048FFFF;
                16'h3494 : rd_rsp_data <= 32'hEBF40004;
                16'h34A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h34A4 : rd_rsp_data <= 32'hEBF40004;
                16'h34B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h34B4 : rd_rsp_data <= 32'hEBF40004;
                16'h34C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h34C4 : rd_rsp_data <= 32'hEBF40004;
                16'h34D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h34D4 : rd_rsp_data <= 32'hEBF40004;
                16'h34E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h34E4 : rd_rsp_data <= 32'hEBF40004;
                16'h34F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h34F4 : rd_rsp_data <= 32'hEBF40004;
                16'h3504 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3508 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h350C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3510 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3514 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3518 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h351C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3520 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3524 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3528 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h352C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3530 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3534 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3538 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h353C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3540 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3544 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3548 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h354C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3550 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3554 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3558 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h355C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3560 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3564 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3568 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h356C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3570 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3574 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3578 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h357C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3580 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3584 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3588 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h358C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3590 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3594 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3598 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h359C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h35FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3600 : rd_rsp_data <= 32'hFEE002F8;
                16'h3610 : rd_rsp_data <= 32'hFEE002F8;
                16'h3620 : rd_rsp_data <= 32'hFEE002F8;
                16'h3630 : rd_rsp_data <= 32'hFEE002F8;
                16'h3640 : rd_rsp_data <= 32'h0020FFFF;
                16'h3644 : rd_rsp_data <= 32'hEBF40004;
                16'h3650 : rd_rsp_data <= 32'h0028FFFF;
                16'h3654 : rd_rsp_data <= 32'hEBF40004;
                16'h3660 : rd_rsp_data <= 32'h0030FFFF;
                16'h3664 : rd_rsp_data <= 32'hEBF40004;
                16'h3670 : rd_rsp_data <= 32'h0038FFFF;
                16'h3674 : rd_rsp_data <= 32'hEBF40004;
                16'h3680 : rd_rsp_data <= 32'h0040FFFF;
                16'h3684 : rd_rsp_data <= 32'hEBF40004;
                16'h3690 : rd_rsp_data <= 32'h0048FFFF;
                16'h3694 : rd_rsp_data <= 32'hEBF40004;
                16'h36A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h36A4 : rd_rsp_data <= 32'hEBF40004;
                16'h36B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h36B4 : rd_rsp_data <= 32'hEBF40004;
                16'h36C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h36C4 : rd_rsp_data <= 32'hEBF40004;
                16'h36D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h36D4 : rd_rsp_data <= 32'hEBF40004;
                16'h36E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h36E4 : rd_rsp_data <= 32'hEBF40004;
                16'h36F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h36F4 : rd_rsp_data <= 32'hEBF40004;
                16'h3704 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3708 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h370C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3710 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3714 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3718 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h371C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3720 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3724 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3728 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h372C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3730 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3734 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3738 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h373C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3740 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3744 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3748 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h374C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3750 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3754 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3758 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h375C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3760 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3764 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3768 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h376C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3770 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3774 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3778 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h377C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3780 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3784 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3788 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h378C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3790 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3794 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3798 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h379C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h37FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3800 : rd_rsp_data <= 32'hFEE002F8;
                16'h3810 : rd_rsp_data <= 32'hFEE002F8;
                16'h3820 : rd_rsp_data <= 32'hFEE002F8;
                16'h3830 : rd_rsp_data <= 32'hFEE002F8;
                16'h3840 : rd_rsp_data <= 32'h0020FFFF;
                16'h3844 : rd_rsp_data <= 32'hEBF40004;
                16'h3850 : rd_rsp_data <= 32'h0028FFFF;
                16'h3854 : rd_rsp_data <= 32'hEBF40004;
                16'h3860 : rd_rsp_data <= 32'h0030FFFF;
                16'h3864 : rd_rsp_data <= 32'hEBF40004;
                16'h3870 : rd_rsp_data <= 32'h0038FFFF;
                16'h3874 : rd_rsp_data <= 32'hEBF40004;
                16'h3880 : rd_rsp_data <= 32'h0040FFFF;
                16'h3884 : rd_rsp_data <= 32'hEBF40004;
                16'h3890 : rd_rsp_data <= 32'h0048FFFF;
                16'h3894 : rd_rsp_data <= 32'hEBF40004;
                16'h38A0 : rd_rsp_data <= 32'h0050FFFF;
                16'h38A4 : rd_rsp_data <= 32'hEBF40004;
                16'h38B0 : rd_rsp_data <= 32'h0058FFFF;
                16'h38B4 : rd_rsp_data <= 32'hEBF40004;
                16'h38C0 : rd_rsp_data <= 32'h0060FFFF;
                16'h38C4 : rd_rsp_data <= 32'hEBF40004;
                16'h38D0 : rd_rsp_data <= 32'h0068FFFF;
                16'h38D4 : rd_rsp_data <= 32'hEBF40004;
                16'h38E0 : rd_rsp_data <= 32'h0070FFFF;
                16'h38E4 : rd_rsp_data <= 32'hEBF40004;
                16'h38F0 : rd_rsp_data <= 32'h0078FFFF;
                16'h38F4 : rd_rsp_data <= 32'hEBF40004;
                16'h3904 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3908 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h390C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3910 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3914 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3918 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h391C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3920 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3924 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3928 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h392C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3930 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3934 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3938 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h393C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3940 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3944 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3948 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h394C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3950 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3954 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3958 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h395C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3960 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3964 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3968 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h396C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3970 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3974 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3978 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h397C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3980 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3984 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3988 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h398C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3990 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3994 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3998 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h399C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39A0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39A4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39A8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39AC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39B0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39B4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39B8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39BC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39C0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39C4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39C8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39CC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39D0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39D4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39D8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39DC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39E0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39E4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39E8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39EC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39F0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39F4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39F8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h39FC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3A00 : rd_rsp_data <= 32'hFEE002F8;
                16'h3A10 : rd_rsp_data <= 32'hFEE002F8;
                16'h3A20 : rd_rsp_data <= 32'hFEE002F8;
                16'h3A30 : rd_rsp_data <= 32'hFEE002F8;
                16'h3A40 : rd_rsp_data <= 32'h0020FFFF;
                16'h3A44 : rd_rsp_data <= 32'hEBF40004;
                16'h3A50 : rd_rsp_data <= 32'h0028FFFF;
                16'h3A54 : rd_rsp_data <= 32'hEBF40004;
                16'h3A60 : rd_rsp_data <= 32'h0030FFFF;
                16'h3A64 : rd_rsp_data <= 32'hEBF40004;
                16'h3A70 : rd_rsp_data <= 32'h0038FFFF;
                16'h3A74 : rd_rsp_data <= 32'hEBF40004;
                16'h3A80 : rd_rsp_data <= 32'h0040FFFF;
                16'h3A84 : rd_rsp_data <= 32'hEBF40004;
                16'h3A90 : rd_rsp_data <= 32'h0048FFFF;
                16'h3A94 : rd_rsp_data <= 32'hEBF40004;
                16'h3AA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h3AA4 : rd_rsp_data <= 32'hEBF40004;
                16'h3AB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h3AB4 : rd_rsp_data <= 32'hEBF40004;
                16'h3AC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h3AC4 : rd_rsp_data <= 32'hEBF40004;
                16'h3AD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h3AD4 : rd_rsp_data <= 32'hEBF40004;
                16'h3AE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h3AE4 : rd_rsp_data <= 32'hEBF40004;
                16'h3AF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h3AF4 : rd_rsp_data <= 32'hEBF40004;
                16'h3B04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3B9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3BFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3C00 : rd_rsp_data <= 32'hFEE002F8;
                16'h3C10 : rd_rsp_data <= 32'hFEE002F8;
                16'h3C20 : rd_rsp_data <= 32'hFEE002F8;
                16'h3C30 : rd_rsp_data <= 32'hFEE002F8;
                16'h3C40 : rd_rsp_data <= 32'h0020FFFF;
                16'h3C44 : rd_rsp_data <= 32'hEBF40004;
                16'h3C50 : rd_rsp_data <= 32'h0028FFFF;
                16'h3C54 : rd_rsp_data <= 32'hEBF40004;
                16'h3C60 : rd_rsp_data <= 32'h0030FFFF;
                16'h3C64 : rd_rsp_data <= 32'hEBF40004;
                16'h3C70 : rd_rsp_data <= 32'h0038FFFF;
                16'h3C74 : rd_rsp_data <= 32'hEBF40004;
                16'h3C80 : rd_rsp_data <= 32'h0040FFFF;
                16'h3C84 : rd_rsp_data <= 32'hEBF40004;
                16'h3C90 : rd_rsp_data <= 32'h0048FFFF;
                16'h3C94 : rd_rsp_data <= 32'hEBF40004;
                16'h3CA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h3CA4 : rd_rsp_data <= 32'hEBF40004;
                16'h3CB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h3CB4 : rd_rsp_data <= 32'hEBF40004;
                16'h3CC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h3CC4 : rd_rsp_data <= 32'hEBF40004;
                16'h3CD0 : rd_rsp_data <= 32'h0068FFFF;
                16'h3CD4 : rd_rsp_data <= 32'hEBF40004;
                16'h3CE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h3CE4 : rd_rsp_data <= 32'hEBF40004;
                16'h3CF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h3CF4 : rd_rsp_data <= 32'hEBF40004;
                16'h3D04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3D9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3DFC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3E00 : rd_rsp_data <= 32'hFEE002F8;
                16'h3E10 : rd_rsp_data <= 32'hFEE002F8;
                16'h3E20 : rd_rsp_data <= 32'hFEE002F8;
                16'h3E30 : rd_rsp_data <= 32'hFEE002F8;
                16'h3E40 : rd_rsp_data <= 32'h0020FFFF;
                16'h3E44 : rd_rsp_data <= 32'hEBF40004;
                16'h3E50 : rd_rsp_data <= 32'h0028FFFF;
                16'h3E54 : rd_rsp_data <= 32'hEBF40004;
                16'h3E60 : rd_rsp_data <= 32'h0030FFFF;
                16'h3E64 : rd_rsp_data <= 32'hEBF40004;
                16'h3E70 : rd_rsp_data <= 32'h0038FFFF;
                16'h3E74 : rd_rsp_data <= 32'hEBF40004;
                16'h3E80 : rd_rsp_data <= 32'h0040FFFF;
                16'h3E84 : rd_rsp_data <= 32'hEBF40004;
                16'h3E90 : rd_rsp_data <= 32'h0048FFFF;
                16'h3E94 : rd_rsp_data <= 32'hEBF40004;
                16'h3EA0 : rd_rsp_data <= 32'h0050FFFF;
                16'h3EA4 : rd_rsp_data <= 32'hEBF40004;
                16'h3EB0 : rd_rsp_data <= 32'h0058FFFF;
                16'h3EB4 : rd_rsp_data <= 32'hEBF40004;
                16'h3EC0 : rd_rsp_data <= 32'h0060FFFF;
                16'h3EC4 : rd_rsp_data <= 32'hEBF40004;
                16'h3ED0 : rd_rsp_data <= 32'h0068FFFF;
                16'h3ED4 : rd_rsp_data <= 32'hEBF40004;
                16'h3EE0 : rd_rsp_data <= 32'h0070FFFF;
                16'h3EE4 : rd_rsp_data <= 32'hEBF40004;
                16'h3EF0 : rd_rsp_data <= 32'h0078FFFF;
                16'h3EF4 : rd_rsp_data <= 32'hEBF40004;
                16'h3F04 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F08 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F0C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F10 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F14 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F18 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F1C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F20 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F24 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F28 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F2C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F30 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F34 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F38 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F3C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F40 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F44 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F48 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F4C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F50 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F54 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F58 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F5C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F60 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F64 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F68 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F6C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F70 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F74 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F78 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F7C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F80 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F84 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F88 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F8C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F90 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F94 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F98 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3F9C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FA0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FA4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FA8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FAC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FB0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FB4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FB8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FBC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FC0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FC4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FC8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FCC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FD0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FD4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FD8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FDC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FE0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FE4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FE8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FEC : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FF0 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FF4 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FF8 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h3FFC : rd_rsp_data <= 32'hFFFFFFFF;
                default: rd_rsp_data <= 32'h00000000;
            endcase
        end else if (dwr_valid) begin
            case (({dwr_addr[31:24], dwr_addr[23:16], dwr_addr[15:08], dwr_addr[07:00]} - (base_address_register & 32'hFFFFFFF0)) & 32'hFFFF)
                //Dont be scared
            endcase
        end else begin
            rd_rsp_data <= 32'h00000000;
        end
    end
            
endmodule
